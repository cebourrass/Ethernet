-- nios_system.vhd

-- Generated using ACDS version 13.0 156 at 2013.10.09.16:22:30

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity nios_system is
	port (
		clk_clk                                      : in  std_logic                     := '0';             --                         clk.clk
		reset_reset_n                                : in  std_logic                     := '0';             --                       reset.reset_n
		pio_0_external_connection_export             : out std_logic;                                        --   pio_0_external_connection.export
		av_status_reg_0_conduit_end_udp_send         : out std_logic;                                        -- av_status_reg_0_conduit_end.udp_send
		av_status_reg_0_conduit_end_status_reg0_o    : out std_logic_vector(31 downto 0);                    --                            .status_reg0_o
		av_status_reg_0_conduit_end_status_reg1_o    : out std_logic_vector(31 downto 0);                    --                            .status_reg1_o
		av_status_reg_0_conduit_end_status_reg2_o    : out std_logic_vector(31 downto 0);                    --                            .status_reg2_o
		av_status_reg_0_conduit_end_status_reg3_o    : out std_logic_vector(31 downto 0);                    --                            .status_reg3_o
		av_status_reg_0_conduit_end_status_reg4_o    : out std_logic_vector(31 downto 0);                    --                            .status_reg4_o
		av_status_reg_0_conduit_end_status_reg5_o    : out std_logic_vector(31 downto 0);                    --                            .status_reg5_o
		av_status_reg_0_conduit_end_status_reg7_o    : out std_logic_vector(31 downto 0);                    --                            .status_reg7_o
		av_status_reg_0_conduit_end_status_reg6_o    : out std_logic_vector(31 downto 0);                    --                            .status_reg6_o
		av_eth_config_0_conduit_end_local_port_o     : out std_logic_vector(15 downto 0);                    -- av_eth_config_0_conduit_end.local_port_o
		av_eth_config_0_conduit_end_remote_port_o    : out std_logic_vector(15 downto 0);                    --                            .remote_port_o
		av_eth_config_0_conduit_end_local_IP_o       : out std_logic_vector(31 downto 0);                    --                            .local_IP_o
		av_eth_config_0_conduit_end_remote_IP_o      : out std_logic_vector(31 downto 0);                    --                            .remote_IP_o
		av_eth_config_0_conduit_end_local_MAC_LSB_o  : out std_logic_vector(31 downto 0);                    --                            .local_MAC_LSB_o
		av_eth_config_0_conduit_end_local_MAC_MSB_o  : out std_logic_vector(31 downto 0);                    --                            .local_MAC_MSB_o
		av_eth_config_0_conduit_end_remote_MAC_LSB_o : out std_logic_vector(31 downto 0);                    --                            .remote_MAC_LSB_o
		av_eth_config_0_conduit_end_checksum_o       : out std_logic_vector(15 downto 0);                    --                            .checksum_o
		av_eth_config_0_conduit_end_remote_MAC_MSB_o : out std_logic_vector(31 downto 0);                    --                            .remote_MAC_MSB_o
		av_config_reg_0_conduit_end_reg_0            : in  std_logic_vector(31 downto 0) := (others => '0'); -- av_config_reg_0_conduit_end.reg_0
		av_config_reg_0_conduit_end_reg_1            : in  std_logic_vector(31 downto 0) := (others => '0'); --                            .reg_1
		av_config_reg_0_conduit_end_reg_2            : in  std_logic_vector(31 downto 0) := (others => '0'); --                            .reg_2
		av_config_reg_0_conduit_end_reg_3            : in  std_logic_vector(31 downto 0) := (others => '0'); --                            .reg_3
		av_config_reg_0_conduit_end_reg_4            : in  std_logic_vector(31 downto 0) := (others => '0'); --                            .reg_4
		av_config_reg_0_conduit_end_reg_5            : in  std_logic_vector(31 downto 0) := (others => '0'); --                            .reg_5
		av_config_reg_0_conduit_end_reg_6            : in  std_logic_vector(31 downto 0) := (others => '0'); --                            .reg_6
		av_config_reg_0_conduit_end_reg_7            : in  std_logic_vector(31 downto 0) := (others => '0'); --                            .reg_7
		av_config_reg_0_conduit_end_udp_data_valid   : in  std_logic                     := '0';             --                            .udp_data_valid
		av_sendpacket_0_conduit_end_checksum_o       : out std_logic_vector(15 downto 0);                    -- av_sendpacket_0_conduit_end.checksum_o
		av_sendpacket_0_conduit_end_local_port_o     : out std_logic_vector(15 downto 0);                    --                            .local_port_o
		av_sendpacket_0_conduit_end_remote_port_o    : out std_logic_vector(15 downto 0);                    --                            .remote_port_o
		av_sendpacket_0_conduit_end_remote_MAC_MSB_o : out std_logic_vector(31 downto 0);                    --                            .remote_MAC_MSB_o
		av_sendpacket_0_conduit_end_remote_MAC_LSB_o : out std_logic_vector(31 downto 0);                    --                            .remote_MAC_LSB_o
		av_sendpacket_0_conduit_end_udp_sendpacket   : out std_logic;                                        --                            .udp_sendpacket
		av_sendpacket_0_conduit_end_length_o         : out std_logic_vector(15 downto 0);                    --                            .length_o
		av_sendpacket_0_conduit_end_remote_IP_o      : out std_logic_vector(31 downto 0)                     --                            .remote_IP_o
	);
end entity nios_system;

architecture rtl of nios_system is
	component nios_system_onchip_memory2_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X'              -- reset
		);
	end component nios_system_onchip_memory2_0;

	component nios_system_nios2_qsys_0 is
		port (
			clk                                   : in  std_logic                     := 'X';             -- clk
			reset_n                               : in  std_logic                     := 'X';             -- reset_n
			d_address                             : out std_logic_vector(19 downto 0);                    -- address
			d_byteenable                          : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                                : out std_logic;                                        -- read
			d_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_write                               : out std_logic;                                        -- write
			d_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_debug_module_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                             : out std_logic_vector(19 downto 0);                    -- address
			i_read                                : out std_logic;                                        -- read
			i_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			jtag_debug_module_resetrequest        : out std_logic;                                        -- reset
			jtag_debug_module_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			jtag_debug_module_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			jtag_debug_module_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			jtag_debug_module_read                : in  std_logic                     := 'X';             -- read
			jtag_debug_module_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			jtag_debug_module_waitrequest         : out std_logic;                                        -- waitrequest
			jtag_debug_module_write               : in  std_logic                     := 'X';             -- write
			jtag_debug_module_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			no_ci_readra                          : out std_logic                                         -- readra
		);
	end component nios_system_nios2_qsys_0;

	component nios_system_jtag_uart_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component nios_system_jtag_uart_0;

	component nios_system_sysid_qsys_0 is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component nios_system_sysid_qsys_0;

	component nios_system_timer_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component nios_system_timer_0;

	component nios_system_pio_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic                                         -- export
		);
	end component nios_system_pio_0;

	component av_status_reg is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			address       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			write         : in  std_logic                     := 'X';             -- write
			read          : in  std_logic                     := 'X';             -- read
			writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			udp_send      : out std_logic;                                        -- export
			status_reg0_o : out std_logic_vector(31 downto 0);                    -- export
			status_reg1_o : out std_logic_vector(31 downto 0);                    -- export
			status_reg2_o : out std_logic_vector(31 downto 0);                    -- export
			status_reg3_o : out std_logic_vector(31 downto 0);                    -- export
			status_reg4_o : out std_logic_vector(31 downto 0);                    -- export
			status_reg5_o : out std_logic_vector(31 downto 0);                    -- export
			status_reg7_o : out std_logic_vector(31 downto 0);                    -- export
			status_reg6_o : out std_logic_vector(31 downto 0)                     -- export
		);
	end component av_status_reg;

	component av_eth_config is
		port (
			clk              : in  std_logic                     := 'X';             -- clk
			reset_n          : in  std_logic                     := 'X';             -- reset_n
			write            : in  std_logic                     := 'X';             -- write
			read             : in  std_logic                     := 'X';             -- read
			writedata        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			address          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			readdata         : out std_logic_vector(31 downto 0);                    -- readdata
			local_port_o     : out std_logic_vector(15 downto 0);                    -- export
			remote_port_o    : out std_logic_vector(15 downto 0);                    -- export
			local_IP_o       : out std_logic_vector(31 downto 0);                    -- export
			remote_IP_o      : out std_logic_vector(31 downto 0);                    -- export
			local_MAC_LSB_o  : out std_logic_vector(31 downto 0);                    -- export
			local_MAC_MSB_o  : out std_logic_vector(31 downto 0);                    -- export
			remote_MAC_LSB_o : out std_logic_vector(31 downto 0);                    -- export
			checksum_o       : out std_logic_vector(15 downto 0);                    -- export
			remote_MAC_MSB_o : out std_logic_vector(31 downto 0)                     -- export
		);
	end component av_eth_config;

	component av_config_reg is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			reset_n        : in  std_logic                     := 'X';             -- reset_n
			address        : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			write          : in  std_logic                     := 'X';             -- write
			read           : in  std_logic                     := 'X';             -- read
			writedata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			reg_0          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- export
			reg_1          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- export
			reg_2          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- export
			reg_3          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- export
			reg_4          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- export
			reg_5          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- export
			reg_6          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- export
			reg_7          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- export
			udp_data_valid : in  std_logic                     := 'X';             -- export
			av_irq         : out std_logic                                         -- irq
		);
	end component av_config_reg;

	component av_sendpacket is
		port (
			clk              : in  std_logic                     := 'X';             -- clk
			reset_n          : in  std_logic                     := 'X';             -- reset_n
			address          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			write            : in  std_logic                     := 'X';             -- write
			read             : in  std_logic                     := 'X';             -- read
			writedata        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata         : out std_logic_vector(31 downto 0);                    -- readdata
			checksum_o       : out std_logic_vector(15 downto 0);                    -- export
			local_port_o     : out std_logic_vector(15 downto 0);                    -- export
			remote_port_o    : out std_logic_vector(15 downto 0);                    -- export
			remote_MAC_MSB_o : out std_logic_vector(31 downto 0);                    -- export
			remote_MAC_LSB_o : out std_logic_vector(31 downto 0);                    -- export
			udp_sendpacket   : out std_logic;                                        -- export
			length_o         : out std_logic_vector(15 downto 0);                    -- export
			remote_IP_o      : out std_logic_vector(31 downto 0)                     -- export
		);
	end component av_sendpacket;

	component altera_merlin_master_agent is
		generic (
			PKT_PROTECTION_H          : integer := 80;
			PKT_PROTECTION_L          : integer := 80;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_BURSTWRAP_H           : integer := 79;
			PKT_BURSTWRAP_L           : integer := 77;
			PKT_BURST_SIZE_H          : integer := 86;
			PKT_BURST_SIZE_L          : integer := 84;
			PKT_BURST_TYPE_H          : integer := 94;
			PKT_BURST_TYPE_L          : integer := 93;
			PKT_BYTE_CNT_H            : integer := 76;
			PKT_BYTE_CNT_L            : integer := 74;
			PKT_ADDR_H                : integer := 73;
			PKT_ADDR_L                : integer := 42;
			PKT_TRANS_COMPRESSED_READ : integer := 41;
			PKT_TRANS_POSTED          : integer := 40;
			PKT_TRANS_WRITE           : integer := 39;
			PKT_TRANS_READ            : integer := 38;
			PKT_TRANS_LOCK            : integer := 82;
			PKT_TRANS_EXCLUSIVE       : integer := 83;
			PKT_DATA_H                : integer := 37;
			PKT_DATA_L                : integer := 6;
			PKT_BYTEEN_H              : integer := 5;
			PKT_BYTEEN_L              : integer := 2;
			PKT_SRC_ID_H              : integer := 1;
			PKT_SRC_ID_L              : integer := 1;
			PKT_DEST_ID_H             : integer := 0;
			PKT_DEST_ID_L             : integer := 0;
			PKT_THREAD_ID_H           : integer := 88;
			PKT_THREAD_ID_L           : integer := 87;
			PKT_CACHE_H               : integer := 92;
			PKT_CACHE_L               : integer := 89;
			PKT_DATA_SIDEBAND_H       : integer := 105;
			PKT_DATA_SIDEBAND_L       : integer := 98;
			PKT_QOS_H                 : integer := 109;
			PKT_QOS_L                 : integer := 106;
			PKT_ADDR_SIDEBAND_H       : integer := 97;
			PKT_ADDR_SIDEBAND_L       : integer := 93;
			PKT_RESPONSE_STATUS_H     : integer := 111;
			PKT_RESPONSE_STATUS_L     : integer := 110;
			ST_DATA_W                 : integer := 112;
			ST_CHANNEL_W              : integer := 1;
			AV_BURSTCOUNT_W           : integer := 3;
			SUPPRESS_0_BYTEEN_RSP     : integer := 1;
			ID                        : integer := 1;
			BURSTWRAP_VALUE           : integer := 4;
			CACHE_VALUE               : integer := 0;
			SECURE_ACCESS_BIT         : integer := 1;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			av_address              : in  std_logic_vector(19 downto 0) := (others => 'X'); -- address
			av_write                : in  std_logic                     := 'X';             -- write
			av_read                 : in  std_logic                     := 'X';             -- read
			av_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			av_waitrequest          : out std_logic;                                        -- waitrequest
			av_readdatavalid        : out std_logic;                                        -- readdatavalid
			av_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			av_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_lock                 : in  std_logic                     := 'X';             -- lock
			cp_valid                : out std_logic;                                        -- valid
			cp_data                 : out std_logic_vector(94 downto 0);                    -- data
			cp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_endofpacket          : out std_logic;                                        -- endofpacket
			cp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : in  std_logic                     := 'X';             -- valid
			rp_data                 : in  std_logic_vector(94 downto 0) := (others => 'X'); -- data
			rp_channel              : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			rp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			rp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			rp_ready                : out std_logic;                                        -- ready
			av_response             : out std_logic_vector(1 downto 0);                     -- response
			av_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid   : out std_logic                                         -- writeresponsevalid
		);
	end component altera_merlin_master_agent;

	component altera_merlin_slave_agent is
		generic (
			PKT_DATA_H                : integer := 31;
			PKT_DATA_L                : integer := 0;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_SYMBOL_W              : integer := 8;
			PKT_BYTEEN_H              : integer := 71;
			PKT_BYTEEN_L              : integer := 68;
			PKT_ADDR_H                : integer := 63;
			PKT_ADDR_L                : integer := 32;
			PKT_TRANS_COMPRESSED_READ : integer := 67;
			PKT_TRANS_POSTED          : integer := 66;
			PKT_TRANS_WRITE           : integer := 65;
			PKT_TRANS_READ            : integer := 64;
			PKT_TRANS_LOCK            : integer := 87;
			PKT_SRC_ID_H              : integer := 74;
			PKT_SRC_ID_L              : integer := 72;
			PKT_DEST_ID_H             : integer := 77;
			PKT_DEST_ID_L             : integer := 75;
			PKT_BURSTWRAP_H           : integer := 85;
			PKT_BURSTWRAP_L           : integer := 82;
			PKT_BYTE_CNT_H            : integer := 81;
			PKT_BYTE_CNT_L            : integer := 78;
			PKT_PROTECTION_H          : integer := 86;
			PKT_PROTECTION_L          : integer := 86;
			PKT_RESPONSE_STATUS_H     : integer := 89;
			PKT_RESPONSE_STATUS_L     : integer := 88;
			PKT_BURST_SIZE_H          : integer := 92;
			PKT_BURST_SIZE_L          : integer := 90;
			ST_CHANNEL_W              : integer := 8;
			ST_DATA_W                 : integer := 93;
			AVS_BURSTCOUNT_W          : integer := 4;
			SUPPRESS_0_BYTEEN_CMD     : integer := 1;
			PREVENT_FIFO_OVERFLOW     : integer := 0;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			m0_address              : out std_logic_vector(19 downto 0);                    -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess          : out std_logic;                                        -- debugaccess
			m0_lock                 : out std_logic;                                        -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                        -- read
			m0_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			m0_write                : out std_logic;                                        -- write
			rp_endofpacket          : out std_logic;                                        -- endofpacket
			rp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : out std_logic;                                        -- valid
			rp_data                 : out std_logic_vector(94 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_ready                : out std_logic;                                        -- ready
			cp_valid                : in  std_logic                     := 'X';             -- valid
			cp_data                 : in  std_logic_vector(94 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                        -- ready
			rf_sink_valid           : in  std_logic                     := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(95 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                     := 'X';             -- ready
			rf_source_valid         : out std_logic;                                        -- valid
			rf_source_startofpacket : out std_logic;                                        -- startofpacket
			rf_source_endofpacket   : out std_logic;                                        -- endofpacket
			rf_source_data          : out std_logic_vector(95 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                        -- ready
			rdata_fifo_sink_valid   : in  std_logic                     := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(33 downto 0) := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                     := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                        -- valid
			rdata_fifo_src_data     : out std_logic_vector(33 downto 0);                    -- data
			m0_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			m0_writeresponserequest : out std_logic;                                        -- writeresponserequest
			m0_writeresponsevalid   : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component altera_merlin_slave_agent;

	component altera_avalon_sc_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			in_data           : in  std_logic_vector(95 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                     := 'X';             -- valid
			in_ready          : out std_logic;                                        -- ready
			in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			out_data          : out std_logic_vector(95 downto 0);                    -- data
			out_valid         : out std_logic;                                        -- valid
			out_ready         : in  std_logic                     := 'X';             -- ready
			out_startofpacket : out std_logic;                                        -- startofpacket
			out_endofpacket   : out std_logic;                                        -- endofpacket
			csr_address       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			csr_read          : in  std_logic                     := 'X';             -- read
			csr_write         : in  std_logic                     := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                        -- data
			almost_empty_data : out std_logic;                                        -- data
			in_empty          : in  std_logic                     := 'X';             -- empty
			out_empty         : out std_logic;                                        -- empty
			in_error          : in  std_logic                     := 'X';             -- error
			out_error         : out std_logic;                                        -- error
			in_channel        : in  std_logic                     := 'X';             -- channel
			out_channel       : out std_logic                                         -- channel
		);
	end component altera_avalon_sc_fifo;

	component nios_system_addr_router is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(94 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(94 downto 0);                    -- data
			src_channel        : out std_logic_vector(9 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component nios_system_addr_router;

	component nios_system_addr_router_001 is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(94 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(94 downto 0);                    -- data
			src_channel        : out std_logic_vector(9 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component nios_system_addr_router_001;

	component nios_system_id_router is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(94 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(94 downto 0);                    -- data
			src_channel        : out std_logic_vector(9 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component nios_system_id_router;

	component nios_system_id_router_002 is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(94 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(94 downto 0);                    -- data
			src_channel        : out std_logic_vector(9 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component nios_system_id_router_002;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS        : integer := 6;
			OUTPUT_RESET_SYNC_EDGES : string  := "deassert";
			SYNC_DEPTH              : integer := 2
		);
		port (
			reset_in0  : in  std_logic := 'X'; -- reset
			clk        : in  std_logic := 'X'; -- clk
			reset_out  : out std_logic;        -- reset
			reset_in1  : in  std_logic := 'X'; -- reset
			reset_in2  : in  std_logic := 'X'; -- reset
			reset_in3  : in  std_logic := 'X'; -- reset
			reset_in4  : in  std_logic := 'X'; -- reset
			reset_in5  : in  std_logic := 'X'; -- reset
			reset_in6  : in  std_logic := 'X'; -- reset
			reset_in7  : in  std_logic := 'X'; -- reset
			reset_in8  : in  std_logic := 'X'; -- reset
			reset_in9  : in  std_logic := 'X'; -- reset
			reset_in10 : in  std_logic := 'X'; -- reset
			reset_in11 : in  std_logic := 'X'; -- reset
			reset_in12 : in  std_logic := 'X'; -- reset
			reset_in13 : in  std_logic := 'X'; -- reset
			reset_in14 : in  std_logic := 'X'; -- reset
			reset_in15 : in  std_logic := 'X'  -- reset
		);
	end component altera_reset_controller;

	component nios_system_cmd_xbar_demux is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			sink_ready         : out std_logic;                                        -- ready
			sink_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(94 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- valid
			src0_ready         : in  std_logic                     := 'X';             -- ready
			src0_valid         : out std_logic;                                        -- valid
			src0_data          : out std_logic_vector(94 downto 0);                    -- data
			src0_channel       : out std_logic_vector(9 downto 0);                     -- channel
			src0_startofpacket : out std_logic;                                        -- startofpacket
			src0_endofpacket   : out std_logic;                                        -- endofpacket
			src1_ready         : in  std_logic                     := 'X';             -- ready
			src1_valid         : out std_logic;                                        -- valid
			src1_data          : out std_logic_vector(94 downto 0);                    -- data
			src1_channel       : out std_logic_vector(9 downto 0);                     -- channel
			src1_startofpacket : out std_logic;                                        -- startofpacket
			src1_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component nios_system_cmd_xbar_demux;

	component nios_system_cmd_xbar_demux_001 is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			sink_ready         : out std_logic;                                        -- ready
			sink_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(94 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- valid
			src0_ready         : in  std_logic                     := 'X';             -- ready
			src0_valid         : out std_logic;                                        -- valid
			src0_data          : out std_logic_vector(94 downto 0);                    -- data
			src0_channel       : out std_logic_vector(9 downto 0);                     -- channel
			src0_startofpacket : out std_logic;                                        -- startofpacket
			src0_endofpacket   : out std_logic;                                        -- endofpacket
			src1_ready         : in  std_logic                     := 'X';             -- ready
			src1_valid         : out std_logic;                                        -- valid
			src1_data          : out std_logic_vector(94 downto 0);                    -- data
			src1_channel       : out std_logic_vector(9 downto 0);                     -- channel
			src1_startofpacket : out std_logic;                                        -- startofpacket
			src1_endofpacket   : out std_logic;                                        -- endofpacket
			src2_ready         : in  std_logic                     := 'X';             -- ready
			src2_valid         : out std_logic;                                        -- valid
			src2_data          : out std_logic_vector(94 downto 0);                    -- data
			src2_channel       : out std_logic_vector(9 downto 0);                     -- channel
			src2_startofpacket : out std_logic;                                        -- startofpacket
			src2_endofpacket   : out std_logic;                                        -- endofpacket
			src3_ready         : in  std_logic                     := 'X';             -- ready
			src3_valid         : out std_logic;                                        -- valid
			src3_data          : out std_logic_vector(94 downto 0);                    -- data
			src3_channel       : out std_logic_vector(9 downto 0);                     -- channel
			src3_startofpacket : out std_logic;                                        -- startofpacket
			src3_endofpacket   : out std_logic;                                        -- endofpacket
			src4_ready         : in  std_logic                     := 'X';             -- ready
			src4_valid         : out std_logic;                                        -- valid
			src4_data          : out std_logic_vector(94 downto 0);                    -- data
			src4_channel       : out std_logic_vector(9 downto 0);                     -- channel
			src4_startofpacket : out std_logic;                                        -- startofpacket
			src4_endofpacket   : out std_logic;                                        -- endofpacket
			src5_ready         : in  std_logic                     := 'X';             -- ready
			src5_valid         : out std_logic;                                        -- valid
			src5_data          : out std_logic_vector(94 downto 0);                    -- data
			src5_channel       : out std_logic_vector(9 downto 0);                     -- channel
			src5_startofpacket : out std_logic;                                        -- startofpacket
			src5_endofpacket   : out std_logic;                                        -- endofpacket
			src6_ready         : in  std_logic                     := 'X';             -- ready
			src6_valid         : out std_logic;                                        -- valid
			src6_data          : out std_logic_vector(94 downto 0);                    -- data
			src6_channel       : out std_logic_vector(9 downto 0);                     -- channel
			src6_startofpacket : out std_logic;                                        -- startofpacket
			src6_endofpacket   : out std_logic;                                        -- endofpacket
			src7_ready         : in  std_logic                     := 'X';             -- ready
			src7_valid         : out std_logic;                                        -- valid
			src7_data          : out std_logic_vector(94 downto 0);                    -- data
			src7_channel       : out std_logic_vector(9 downto 0);                     -- channel
			src7_startofpacket : out std_logic;                                        -- startofpacket
			src7_endofpacket   : out std_logic;                                        -- endofpacket
			src8_ready         : in  std_logic                     := 'X';             -- ready
			src8_valid         : out std_logic;                                        -- valid
			src8_data          : out std_logic_vector(94 downto 0);                    -- data
			src8_channel       : out std_logic_vector(9 downto 0);                     -- channel
			src8_startofpacket : out std_logic;                                        -- startofpacket
			src8_endofpacket   : out std_logic;                                        -- endofpacket
			src9_ready         : in  std_logic                     := 'X';             -- ready
			src9_valid         : out std_logic;                                        -- valid
			src9_data          : out std_logic_vector(94 downto 0);                    -- data
			src9_channel       : out std_logic_vector(9 downto 0);                     -- channel
			src9_startofpacket : out std_logic;                                        -- startofpacket
			src9_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component nios_system_cmd_xbar_demux_001;

	component nios_system_cmd_xbar_mux is
		port (
			clk                 : in  std_logic                     := 'X';             -- clk
			reset               : in  std_logic                     := 'X';             -- reset
			src_ready           : in  std_logic                     := 'X';             -- ready
			src_valid           : out std_logic;                                        -- valid
			src_data            : out std_logic_vector(94 downto 0);                    -- data
			src_channel         : out std_logic_vector(9 downto 0);                     -- channel
			src_startofpacket   : out std_logic;                                        -- startofpacket
			src_endofpacket     : out std_logic;                                        -- endofpacket
			sink0_ready         : out std_logic;                                        -- ready
			sink0_valid         : in  std_logic                     := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(94 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                        -- ready
			sink1_valid         : in  std_logic                     := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(94 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                     := 'X'              -- endofpacket
		);
	end component nios_system_cmd_xbar_mux;

	component nios_system_rsp_xbar_demux_002 is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			sink_ready         : out std_logic;                                        -- ready
			sink_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(94 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- valid
			src0_ready         : in  std_logic                     := 'X';             -- ready
			src0_valid         : out std_logic;                                        -- valid
			src0_data          : out std_logic_vector(94 downto 0);                    -- data
			src0_channel       : out std_logic_vector(9 downto 0);                     -- channel
			src0_startofpacket : out std_logic;                                        -- startofpacket
			src0_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component nios_system_rsp_xbar_demux_002;

	component nios_system_rsp_xbar_mux is
		port (
			clk                 : in  std_logic                     := 'X';             -- clk
			reset               : in  std_logic                     := 'X';             -- reset
			src_ready           : in  std_logic                     := 'X';             -- ready
			src_valid           : out std_logic;                                        -- valid
			src_data            : out std_logic_vector(94 downto 0);                    -- data
			src_channel         : out std_logic_vector(9 downto 0);                     -- channel
			src_startofpacket   : out std_logic;                                        -- startofpacket
			src_endofpacket     : out std_logic;                                        -- endofpacket
			sink0_ready         : out std_logic;                                        -- ready
			sink0_valid         : in  std_logic                     := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(94 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                        -- ready
			sink1_valid         : in  std_logic                     := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(94 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                     := 'X'              -- endofpacket
		);
	end component nios_system_rsp_xbar_mux;

	component nios_system_rsp_xbar_mux_001 is
		port (
			clk                 : in  std_logic                     := 'X';             -- clk
			reset               : in  std_logic                     := 'X';             -- reset
			src_ready           : in  std_logic                     := 'X';             -- ready
			src_valid           : out std_logic;                                        -- valid
			src_data            : out std_logic_vector(94 downto 0);                    -- data
			src_channel         : out std_logic_vector(9 downto 0);                     -- channel
			src_startofpacket   : out std_logic;                                        -- startofpacket
			src_endofpacket     : out std_logic;                                        -- endofpacket
			sink0_ready         : out std_logic;                                        -- ready
			sink0_valid         : in  std_logic                     := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(94 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                        -- ready
			sink1_valid         : in  std_logic                     := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(94 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink2_ready         : out std_logic;                                        -- ready
			sink2_valid         : in  std_logic                     := 'X';             -- valid
			sink2_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink2_data          : in  std_logic_vector(94 downto 0) := (others => 'X'); -- data
			sink2_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink2_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink3_ready         : out std_logic;                                        -- ready
			sink3_valid         : in  std_logic                     := 'X';             -- valid
			sink3_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink3_data          : in  std_logic_vector(94 downto 0) := (others => 'X'); -- data
			sink3_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink3_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink4_ready         : out std_logic;                                        -- ready
			sink4_valid         : in  std_logic                     := 'X';             -- valid
			sink4_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink4_data          : in  std_logic_vector(94 downto 0) := (others => 'X'); -- data
			sink4_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink4_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink5_ready         : out std_logic;                                        -- ready
			sink5_valid         : in  std_logic                     := 'X';             -- valid
			sink5_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink5_data          : in  std_logic_vector(94 downto 0) := (others => 'X'); -- data
			sink5_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink5_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink6_ready         : out std_logic;                                        -- ready
			sink6_valid         : in  std_logic                     := 'X';             -- valid
			sink6_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink6_data          : in  std_logic_vector(94 downto 0) := (others => 'X'); -- data
			sink6_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink6_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink7_ready         : out std_logic;                                        -- ready
			sink7_valid         : in  std_logic                     := 'X';             -- valid
			sink7_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink7_data          : in  std_logic_vector(94 downto 0) := (others => 'X'); -- data
			sink7_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink7_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink8_ready         : out std_logic;                                        -- ready
			sink8_valid         : in  std_logic                     := 'X';             -- valid
			sink8_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink8_data          : in  std_logic_vector(94 downto 0) := (others => 'X'); -- data
			sink8_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink8_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink9_ready         : out std_logic;                                        -- ready
			sink9_valid         : in  std_logic                     := 'X';             -- valid
			sink9_channel       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- channel
			sink9_data          : in  std_logic_vector(94 downto 0) := (others => 'X'); -- data
			sink9_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink9_endofpacket   : in  std_logic                     := 'X'              -- endofpacket
		);
	end component nios_system_rsp_xbar_mux_001;

	component nios_system_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component nios_system_irq_mapper;

	component nios_system_nios2_qsys_0_instruction_master_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(19 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(19 downto 0) := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			av_burstcount            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			av_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_lock                  : in  std_logic                     := 'X';             -- lock
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component nios_system_nios2_qsys_0_instruction_master_translator;

	component nios_system_nios2_qsys_0_data_master_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(19 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(19 downto 0) := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			av_burstcount            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_lock                  : in  std_logic                     := 'X';             -- lock
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component nios_system_nios2_qsys_0_data_master_translator;

	component nios_system_nios2_qsys_0_jtag_debug_module_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(19 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(8 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component nios_system_nios2_qsys_0_jtag_debug_module_translator;

	component nios_system_onchip_memory2_0_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(19 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(15 downto 0);                    -- address
			av_write                 : out std_logic;                                        -- write
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			av_read                  : out std_logic;                                        -- read
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component nios_system_onchip_memory2_0_s1_translator;

	component nios_system_jtag_uart_0_avalon_jtag_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(19 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(0 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_chipselect            : out std_logic;                                        -- chipselect
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component nios_system_jtag_uart_0_avalon_jtag_slave_translator;

	component nios_system_sysid_qsys_0_control_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(19 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(0 downto 0);                     -- address
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component nios_system_sysid_qsys_0_control_slave_translator;

	component nios_system_timer_0_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(19 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(2 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_readdata              : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(15 downto 0);                    -- writedata
			av_chipselect            : out std_logic;                                        -- chipselect
			av_read                  : out std_logic;                                        -- read
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component nios_system_timer_0_s1_translator;

	component nios_system_pio_0_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(19 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(1 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_chipselect            : out std_logic;                                        -- chipselect
			av_read                  : out std_logic;                                        -- read
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component nios_system_pio_0_s1_translator;

	component nios_system_av_status_reg_0_avalon_slave_0_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(19 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(3 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component nios_system_av_status_reg_0_avalon_slave_0_translator;

	signal nios2_qsys_0_instruction_master_waitrequest                                                         : std_logic;                     -- nios2_qsys_0_instruction_master_translator:av_waitrequest -> nios2_qsys_0:i_waitrequest
	signal nios2_qsys_0_instruction_master_address                                                             : std_logic_vector(19 downto 0); -- nios2_qsys_0:i_address -> nios2_qsys_0_instruction_master_translator:av_address
	signal nios2_qsys_0_instruction_master_read                                                                : std_logic;                     -- nios2_qsys_0:i_read -> nios2_qsys_0_instruction_master_translator:av_read
	signal nios2_qsys_0_instruction_master_readdata                                                            : std_logic_vector(31 downto 0); -- nios2_qsys_0_instruction_master_translator:av_readdata -> nios2_qsys_0:i_readdata
	signal nios2_qsys_0_data_master_waitrequest                                                                : std_logic;                     -- nios2_qsys_0_data_master_translator:av_waitrequest -> nios2_qsys_0:d_waitrequest
	signal nios2_qsys_0_data_master_writedata                                                                  : std_logic_vector(31 downto 0); -- nios2_qsys_0:d_writedata -> nios2_qsys_0_data_master_translator:av_writedata
	signal nios2_qsys_0_data_master_address                                                                    : std_logic_vector(19 downto 0); -- nios2_qsys_0:d_address -> nios2_qsys_0_data_master_translator:av_address
	signal nios2_qsys_0_data_master_write                                                                      : std_logic;                     -- nios2_qsys_0:d_write -> nios2_qsys_0_data_master_translator:av_write
	signal nios2_qsys_0_data_master_read                                                                       : std_logic;                     -- nios2_qsys_0:d_read -> nios2_qsys_0_data_master_translator:av_read
	signal nios2_qsys_0_data_master_readdata                                                                   : std_logic_vector(31 downto 0); -- nios2_qsys_0_data_master_translator:av_readdata -> nios2_qsys_0:d_readdata
	signal nios2_qsys_0_data_master_debugaccess                                                                : std_logic;                     -- nios2_qsys_0:jtag_debug_module_debugaccess_to_roms -> nios2_qsys_0_data_master_translator:av_debugaccess
	signal nios2_qsys_0_data_master_byteenable                                                                 : std_logic_vector(3 downto 0);  -- nios2_qsys_0:d_byteenable -> nios2_qsys_0_data_master_translator:av_byteenable
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest                           : std_logic;                     -- nios2_qsys_0:jtag_debug_module_waitrequest -> nios2_qsys_0_jtag_debug_module_translator:av_waitrequest
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata                             : std_logic_vector(31 downto 0); -- nios2_qsys_0_jtag_debug_module_translator:av_writedata -> nios2_qsys_0:jtag_debug_module_writedata
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_address                               : std_logic_vector(8 downto 0);  -- nios2_qsys_0_jtag_debug_module_translator:av_address -> nios2_qsys_0:jtag_debug_module_address
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_write                                 : std_logic;                     -- nios2_qsys_0_jtag_debug_module_translator:av_write -> nios2_qsys_0:jtag_debug_module_write
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_read                                  : std_logic;                     -- nios2_qsys_0_jtag_debug_module_translator:av_read -> nios2_qsys_0:jtag_debug_module_read
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata                              : std_logic_vector(31 downto 0); -- nios2_qsys_0:jtag_debug_module_readdata -> nios2_qsys_0_jtag_debug_module_translator:av_readdata
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess                           : std_logic;                     -- nios2_qsys_0_jtag_debug_module_translator:av_debugaccess -> nios2_qsys_0:jtag_debug_module_debugaccess
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable                            : std_logic_vector(3 downto 0);  -- nios2_qsys_0_jtag_debug_module_translator:av_byteenable -> nios2_qsys_0:jtag_debug_module_byteenable
	signal onchip_memory2_0_s1_translator_avalon_anti_slave_0_writedata                                        : std_logic_vector(31 downto 0); -- onchip_memory2_0_s1_translator:av_writedata -> onchip_memory2_0:writedata
	signal onchip_memory2_0_s1_translator_avalon_anti_slave_0_address                                          : std_logic_vector(15 downto 0); -- onchip_memory2_0_s1_translator:av_address -> onchip_memory2_0:address
	signal onchip_memory2_0_s1_translator_avalon_anti_slave_0_chipselect                                       : std_logic;                     -- onchip_memory2_0_s1_translator:av_chipselect -> onchip_memory2_0:chipselect
	signal onchip_memory2_0_s1_translator_avalon_anti_slave_0_clken                                            : std_logic;                     -- onchip_memory2_0_s1_translator:av_clken -> onchip_memory2_0:clken
	signal onchip_memory2_0_s1_translator_avalon_anti_slave_0_write                                            : std_logic;                     -- onchip_memory2_0_s1_translator:av_write -> onchip_memory2_0:write
	signal onchip_memory2_0_s1_translator_avalon_anti_slave_0_readdata                                         : std_logic_vector(31 downto 0); -- onchip_memory2_0:readdata -> onchip_memory2_0_s1_translator:av_readdata
	signal onchip_memory2_0_s1_translator_avalon_anti_slave_0_byteenable                                       : std_logic_vector(3 downto 0);  -- onchip_memory2_0_s1_translator:av_byteenable -> onchip_memory2_0:byteenable
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest                            : std_logic;                     -- jtag_uart_0:av_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator:av_waitrequest
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata                              : std_logic_vector(31 downto 0); -- jtag_uart_0_avalon_jtag_slave_translator:av_writedata -> jtag_uart_0:av_writedata
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address                                : std_logic_vector(0 downto 0);  -- jtag_uart_0_avalon_jtag_slave_translator:av_address -> jtag_uart_0:av_address
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect                             : std_logic;                     -- jtag_uart_0_avalon_jtag_slave_translator:av_chipselect -> jtag_uart_0:av_chipselect
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write                                  : std_logic;                     -- jtag_uart_0_avalon_jtag_slave_translator:av_write -> jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write:in
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read                                   : std_logic;                     -- jtag_uart_0_avalon_jtag_slave_translator:av_read -> jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read:in
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata                               : std_logic_vector(31 downto 0); -- jtag_uart_0:av_readdata -> jtag_uart_0_avalon_jtag_slave_translator:av_readdata
	signal sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_address                                   : std_logic_vector(0 downto 0);  -- sysid_qsys_0_control_slave_translator:av_address -> sysid_qsys_0:address
	signal sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_readdata                                  : std_logic_vector(31 downto 0); -- sysid_qsys_0:readdata -> sysid_qsys_0_control_slave_translator:av_readdata
	signal timer_0_s1_translator_avalon_anti_slave_0_writedata                                                 : std_logic_vector(15 downto 0); -- timer_0_s1_translator:av_writedata -> timer_0:writedata
	signal timer_0_s1_translator_avalon_anti_slave_0_address                                                   : std_logic_vector(2 downto 0);  -- timer_0_s1_translator:av_address -> timer_0:address
	signal timer_0_s1_translator_avalon_anti_slave_0_chipselect                                                : std_logic;                     -- timer_0_s1_translator:av_chipselect -> timer_0:chipselect
	signal timer_0_s1_translator_avalon_anti_slave_0_write                                                     : std_logic;                     -- timer_0_s1_translator:av_write -> timer_0_s1_translator_avalon_anti_slave_0_write:in
	signal timer_0_s1_translator_avalon_anti_slave_0_readdata                                                  : std_logic_vector(15 downto 0); -- timer_0:readdata -> timer_0_s1_translator:av_readdata
	signal pio_0_s1_translator_avalon_anti_slave_0_writedata                                                   : std_logic_vector(31 downto 0); -- pio_0_s1_translator:av_writedata -> pio_0:writedata
	signal pio_0_s1_translator_avalon_anti_slave_0_address                                                     : std_logic_vector(1 downto 0);  -- pio_0_s1_translator:av_address -> pio_0:address
	signal pio_0_s1_translator_avalon_anti_slave_0_chipselect                                                  : std_logic;                     -- pio_0_s1_translator:av_chipselect -> pio_0:chipselect
	signal pio_0_s1_translator_avalon_anti_slave_0_write                                                       : std_logic;                     -- pio_0_s1_translator:av_write -> pio_0_s1_translator_avalon_anti_slave_0_write:in
	signal pio_0_s1_translator_avalon_anti_slave_0_readdata                                                    : std_logic_vector(31 downto 0); -- pio_0:readdata -> pio_0_s1_translator:av_readdata
	signal av_status_reg_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata                             : std_logic_vector(31 downto 0); -- av_status_reg_0_avalon_slave_0_translator:av_writedata -> av_status_reg_0:writedata
	signal av_status_reg_0_avalon_slave_0_translator_avalon_anti_slave_0_address                               : std_logic_vector(3 downto 0);  -- av_status_reg_0_avalon_slave_0_translator:av_address -> av_status_reg_0:address
	signal av_status_reg_0_avalon_slave_0_translator_avalon_anti_slave_0_write                                 : std_logic;                     -- av_status_reg_0_avalon_slave_0_translator:av_write -> av_status_reg_0:write
	signal av_status_reg_0_avalon_slave_0_translator_avalon_anti_slave_0_read                                  : std_logic;                     -- av_status_reg_0_avalon_slave_0_translator:av_read -> av_status_reg_0:read
	signal av_status_reg_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata                              : std_logic_vector(31 downto 0); -- av_status_reg_0:readdata -> av_status_reg_0_avalon_slave_0_translator:av_readdata
	signal av_eth_config_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata                             : std_logic_vector(31 downto 0); -- av_eth_config_0_avalon_slave_0_translator:av_writedata -> av_eth_config_0:writedata
	signal av_eth_config_0_avalon_slave_0_translator_avalon_anti_slave_0_address                               : std_logic_vector(3 downto 0);  -- av_eth_config_0_avalon_slave_0_translator:av_address -> av_eth_config_0:address
	signal av_eth_config_0_avalon_slave_0_translator_avalon_anti_slave_0_write                                 : std_logic;                     -- av_eth_config_0_avalon_slave_0_translator:av_write -> av_eth_config_0:write
	signal av_eth_config_0_avalon_slave_0_translator_avalon_anti_slave_0_read                                  : std_logic;                     -- av_eth_config_0_avalon_slave_0_translator:av_read -> av_eth_config_0:read
	signal av_eth_config_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata                              : std_logic_vector(31 downto 0); -- av_eth_config_0:readdata -> av_eth_config_0_avalon_slave_0_translator:av_readdata
	signal av_config_reg_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata                             : std_logic_vector(31 downto 0); -- av_config_reg_0_avalon_slave_0_translator:av_writedata -> av_config_reg_0:writedata
	signal av_config_reg_0_avalon_slave_0_translator_avalon_anti_slave_0_address                               : std_logic_vector(3 downto 0);  -- av_config_reg_0_avalon_slave_0_translator:av_address -> av_config_reg_0:address
	signal av_config_reg_0_avalon_slave_0_translator_avalon_anti_slave_0_write                                 : std_logic;                     -- av_config_reg_0_avalon_slave_0_translator:av_write -> av_config_reg_0:write
	signal av_config_reg_0_avalon_slave_0_translator_avalon_anti_slave_0_read                                  : std_logic;                     -- av_config_reg_0_avalon_slave_0_translator:av_read -> av_config_reg_0:read
	signal av_config_reg_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata                              : std_logic_vector(31 downto 0); -- av_config_reg_0:readdata -> av_config_reg_0_avalon_slave_0_translator:av_readdata
	signal av_sendpacket_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata                             : std_logic_vector(31 downto 0); -- av_sendpacket_0_avalon_slave_0_translator:av_writedata -> av_sendpacket_0:writedata
	signal av_sendpacket_0_avalon_slave_0_translator_avalon_anti_slave_0_address                               : std_logic_vector(3 downto 0);  -- av_sendpacket_0_avalon_slave_0_translator:av_address -> av_sendpacket_0:address
	signal av_sendpacket_0_avalon_slave_0_translator_avalon_anti_slave_0_write                                 : std_logic;                     -- av_sendpacket_0_avalon_slave_0_translator:av_write -> av_sendpacket_0:write
	signal av_sendpacket_0_avalon_slave_0_translator_avalon_anti_slave_0_read                                  : std_logic;                     -- av_sendpacket_0_avalon_slave_0_translator:av_read -> av_sendpacket_0:read
	signal av_sendpacket_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata                              : std_logic_vector(31 downto 0); -- av_sendpacket_0:readdata -> av_sendpacket_0_avalon_slave_0_translator:av_readdata
	signal nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_waitrequest                    : std_logic;                     -- nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_qsys_0_instruction_master_translator:uav_waitrequest
	signal nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_burstcount                     : std_logic_vector(2 downto 0);  -- nios2_qsys_0_instruction_master_translator:uav_burstcount -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	signal nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_writedata                      : std_logic_vector(31 downto 0); -- nios2_qsys_0_instruction_master_translator:uav_writedata -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	signal nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_address                        : std_logic_vector(19 downto 0); -- nios2_qsys_0_instruction_master_translator:uav_address -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_address
	signal nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_lock                           : std_logic;                     -- nios2_qsys_0_instruction_master_translator:uav_lock -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	signal nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_write                          : std_logic;                     -- nios2_qsys_0_instruction_master_translator:uav_write -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_write
	signal nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_read                           : std_logic;                     -- nios2_qsys_0_instruction_master_translator:uav_read -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_read
	signal nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdata                       : std_logic_vector(31 downto 0); -- nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_qsys_0_instruction_master_translator:uav_readdata
	signal nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_debugaccess                    : std_logic;                     -- nios2_qsys_0_instruction_master_translator:uav_debugaccess -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	signal nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_byteenable                     : std_logic_vector(3 downto 0);  -- nios2_qsys_0_instruction_master_translator:uav_byteenable -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	signal nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdatavalid                  : std_logic;                     -- nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_qsys_0_instruction_master_translator:uav_readdatavalid
	signal nios2_qsys_0_data_master_translator_avalon_universal_master_0_waitrequest                           : std_logic;                     -- nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_qsys_0_data_master_translator:uav_waitrequest
	signal nios2_qsys_0_data_master_translator_avalon_universal_master_0_burstcount                            : std_logic_vector(2 downto 0);  -- nios2_qsys_0_data_master_translator:uav_burstcount -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	signal nios2_qsys_0_data_master_translator_avalon_universal_master_0_writedata                             : std_logic_vector(31 downto 0); -- nios2_qsys_0_data_master_translator:uav_writedata -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_writedata
	signal nios2_qsys_0_data_master_translator_avalon_universal_master_0_address                               : std_logic_vector(19 downto 0); -- nios2_qsys_0_data_master_translator:uav_address -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_address
	signal nios2_qsys_0_data_master_translator_avalon_universal_master_0_lock                                  : std_logic;                     -- nios2_qsys_0_data_master_translator:uav_lock -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_lock
	signal nios2_qsys_0_data_master_translator_avalon_universal_master_0_write                                 : std_logic;                     -- nios2_qsys_0_data_master_translator:uav_write -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_write
	signal nios2_qsys_0_data_master_translator_avalon_universal_master_0_read                                  : std_logic;                     -- nios2_qsys_0_data_master_translator:uav_read -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_read
	signal nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdata                              : std_logic_vector(31 downto 0); -- nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_qsys_0_data_master_translator:uav_readdata
	signal nios2_qsys_0_data_master_translator_avalon_universal_master_0_debugaccess                           : std_logic;                     -- nios2_qsys_0_data_master_translator:uav_debugaccess -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	signal nios2_qsys_0_data_master_translator_avalon_universal_master_0_byteenable                            : std_logic_vector(3 downto 0);  -- nios2_qsys_0_data_master_translator:uav_byteenable -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	signal nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdatavalid                         : std_logic;                     -- nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_qsys_0_data_master_translator:uav_readdatavalid
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest             : std_logic;                     -- nios2_qsys_0_jtag_debug_module_translator:uav_waitrequest -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount              : std_logic_vector(2 downto 0);  -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> nios2_qsys_0_jtag_debug_module_translator:uav_burstcount
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata               : std_logic_vector(31 downto 0); -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> nios2_qsys_0_jtag_debug_module_translator:uav_writedata
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address                 : std_logic_vector(19 downto 0); -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> nios2_qsys_0_jtag_debug_module_translator:uav_address
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write                   : std_logic;                     -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> nios2_qsys_0_jtag_debug_module_translator:uav_write
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock                    : std_logic;                     -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> nios2_qsys_0_jtag_debug_module_translator:uav_lock
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read                    : std_logic;                     -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> nios2_qsys_0_jtag_debug_module_translator:uav_read
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata                : std_logic_vector(31 downto 0); -- nios2_qsys_0_jtag_debug_module_translator:uav_readdata -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid           : std_logic;                     -- nios2_qsys_0_jtag_debug_module_translator:uav_readdatavalid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess             : std_logic;                     -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> nios2_qsys_0_jtag_debug_module_translator:uav_debugaccess
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable              : std_logic_vector(3 downto 0);  -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> nios2_qsys_0_jtag_debug_module_translator:uav_byteenable
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket      : std_logic;                     -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid            : std_logic;                     -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket    : std_logic;                     -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data             : std_logic_vector(95 downto 0); -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready            : std_logic;                     -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket   : std_logic;                     -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid         : std_logic;                     -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket : std_logic;                     -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data          : std_logic_vector(95 downto 0); -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready         : std_logic;                     -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid       : std_logic;                     -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data        : std_logic_vector(33 downto 0); -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready       : std_logic;                     -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                        : std_logic;                     -- onchip_memory2_0_s1_translator:uav_waitrequest -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                         : std_logic_vector(2 downto 0);  -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> onchip_memory2_0_s1_translator:uav_burstcount
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata                          : std_logic_vector(31 downto 0); -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> onchip_memory2_0_s1_translator:uav_writedata
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_address                            : std_logic_vector(19 downto 0); -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> onchip_memory2_0_s1_translator:uav_address
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_write                              : std_logic;                     -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> onchip_memory2_0_s1_translator:uav_write
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_lock                               : std_logic;                     -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> onchip_memory2_0_s1_translator:uav_lock
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_read                               : std_logic;                     -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> onchip_memory2_0_s1_translator:uav_read
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata                           : std_logic_vector(31 downto 0); -- onchip_memory2_0_s1_translator:uav_readdata -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                      : std_logic;                     -- onchip_memory2_0_s1_translator:uav_readdatavalid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                        : std_logic;                     -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> onchip_memory2_0_s1_translator:uav_debugaccess
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                         : std_logic_vector(3 downto 0);  -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> onchip_memory2_0_s1_translator:uav_byteenable
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                 : std_logic;                     -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                       : std_logic;                     -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket               : std_logic;                     -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data                        : std_logic_vector(95 downto 0); -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                       : std_logic;                     -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket              : std_logic;                     -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                    : std_logic;                     -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket            : std_logic;                     -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                     : std_logic_vector(95 downto 0); -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                    : std_logic;                     -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                  : std_logic;                     -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                   : std_logic_vector(33 downto 0); -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                  : std_logic;                     -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest              : std_logic;                     -- jtag_uart_0_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount               : std_logic_vector(2 downto 0);  -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_0_avalon_jtag_slave_translator:uav_burstcount
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata                : std_logic_vector(31 downto 0); -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_0_avalon_jtag_slave_translator:uav_writedata
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address                  : std_logic_vector(19 downto 0); -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_0_avalon_jtag_slave_translator:uav_address
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write                    : std_logic;                     -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_0_avalon_jtag_slave_translator:uav_write
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock                     : std_logic;                     -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_0_avalon_jtag_slave_translator:uav_lock
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read                     : std_logic;                     -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_0_avalon_jtag_slave_translator:uav_read
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata                 : std_logic_vector(31 downto 0); -- jtag_uart_0_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid            : std_logic;                     -- jtag_uart_0_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess              : std_logic;                     -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_0_avalon_jtag_slave_translator:uav_debugaccess
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable               : std_logic_vector(3 downto 0);  -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_0_avalon_jtag_slave_translator:uav_byteenable
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket       : std_logic;                     -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid             : std_logic;                     -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket     : std_logic;                     -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data              : std_logic_vector(95 downto 0); -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready             : std_logic;                     -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    : std_logic;                     -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid          : std_logic;                     -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket  : std_logic;                     -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data           : std_logic_vector(95 downto 0); -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready          : std_logic;                     -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid        : std_logic;                     -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data         : std_logic_vector(33 downto 0); -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready        : std_logic;                     -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest                 : std_logic;                     -- sysid_qsys_0_control_slave_translator:uav_waitrequest -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount                  : std_logic_vector(2 downto 0);  -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sysid_qsys_0_control_slave_translator:uav_burstcount
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata                   : std_logic_vector(31 downto 0); -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sysid_qsys_0_control_slave_translator:uav_writedata
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_address                     : std_logic_vector(19 downto 0); -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> sysid_qsys_0_control_slave_translator:uav_address
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_write                       : std_logic;                     -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> sysid_qsys_0_control_slave_translator:uav_write
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_lock                        : std_logic;                     -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sysid_qsys_0_control_slave_translator:uav_lock
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_read                        : std_logic;                     -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> sysid_qsys_0_control_slave_translator:uav_read
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata                    : std_logic_vector(31 downto 0); -- sysid_qsys_0_control_slave_translator:uav_readdata -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid               : std_logic;                     -- sysid_qsys_0_control_slave_translator:uav_readdatavalid -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess                 : std_logic;                     -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sysid_qsys_0_control_slave_translator:uav_debugaccess
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable                  : std_logic_vector(3 downto 0);  -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sysid_qsys_0_control_slave_translator:uav_byteenable
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket          : std_logic;                     -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid                : std_logic;                     -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket        : std_logic;                     -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data                 : std_logic_vector(95 downto 0); -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready                : std_logic;                     -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket       : std_logic;                     -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid             : std_logic;                     -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket     : std_logic;                     -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data              : std_logic_vector(95 downto 0); -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready             : std_logic;                     -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid           : std_logic;                     -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data            : std_logic_vector(33 downto 0); -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready           : std_logic;                     -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                 : std_logic;                     -- timer_0_s1_translator:uav_waitrequest -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                  : std_logic_vector(2 downto 0);  -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_0_s1_translator:uav_burstcount
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                   : std_logic_vector(31 downto 0); -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_0_s1_translator:uav_writedata
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address                                     : std_logic_vector(19 downto 0); -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_0_s1_translator:uav_address
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write                                       : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_0_s1_translator:uav_write
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock                                        : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_0_s1_translator:uav_lock
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read                                        : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_0_s1_translator:uav_read
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                    : std_logic_vector(31 downto 0); -- timer_0_s1_translator:uav_readdata -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                               : std_logic;                     -- timer_0_s1_translator:uav_readdatavalid -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                 : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_0_s1_translator:uav_debugaccess
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                  : std_logic_vector(3 downto 0);  -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_0_s1_translator:uav_byteenable
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                          : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                        : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                 : std_logic_vector(95 downto 0); -- timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                       : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                             : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                     : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                              : std_logic_vector(95 downto 0); -- timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                             : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                           : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                            : std_logic_vector(33 downto 0); -- timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                           : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal pio_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                   : std_logic;                     -- pio_0_s1_translator:uav_waitrequest -> pio_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal pio_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                    : std_logic_vector(2 downto 0);  -- pio_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_0_s1_translator:uav_burstcount
	signal pio_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                     : std_logic_vector(31 downto 0); -- pio_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_0_s1_translator:uav_writedata
	signal pio_0_s1_translator_avalon_universal_slave_0_agent_m0_address                                       : std_logic_vector(19 downto 0); -- pio_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_0_s1_translator:uav_address
	signal pio_0_s1_translator_avalon_universal_slave_0_agent_m0_write                                         : std_logic;                     -- pio_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_0_s1_translator:uav_write
	signal pio_0_s1_translator_avalon_universal_slave_0_agent_m0_lock                                          : std_logic;                     -- pio_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_0_s1_translator:uav_lock
	signal pio_0_s1_translator_avalon_universal_slave_0_agent_m0_read                                          : std_logic;                     -- pio_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_0_s1_translator:uav_read
	signal pio_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                      : std_logic_vector(31 downto 0); -- pio_0_s1_translator:uav_readdata -> pio_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal pio_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                 : std_logic;                     -- pio_0_s1_translator:uav_readdatavalid -> pio_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal pio_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                   : std_logic;                     -- pio_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_0_s1_translator:uav_debugaccess
	signal pio_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                    : std_logic_vector(3 downto 0);  -- pio_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_0_s1_translator:uav_byteenable
	signal pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                            : std_logic;                     -- pio_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                  : std_logic;                     -- pio_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                          : std_logic;                     -- pio_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                   : std_logic_vector(95 downto 0); -- pio_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                  : std_logic;                     -- pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                         : std_logic;                     -- pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                               : std_logic;                     -- pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                       : std_logic;                     -- pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                : std_logic_vector(95 downto 0); -- pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                               : std_logic;                     -- pio_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                             : std_logic;                     -- pio_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                              : std_logic_vector(33 downto 0); -- pio_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                             : std_logic;                     -- pio_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest             : std_logic;                     -- av_status_reg_0_avalon_slave_0_translator:uav_waitrequest -> av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount              : std_logic_vector(2 downto 0);  -- av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> av_status_reg_0_avalon_slave_0_translator:uav_burstcount
	signal av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata               : std_logic_vector(31 downto 0); -- av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> av_status_reg_0_avalon_slave_0_translator:uav_writedata
	signal av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address                 : std_logic_vector(19 downto 0); -- av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> av_status_reg_0_avalon_slave_0_translator:uav_address
	signal av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write                   : std_logic;                     -- av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> av_status_reg_0_avalon_slave_0_translator:uav_write
	signal av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock                    : std_logic;                     -- av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> av_status_reg_0_avalon_slave_0_translator:uav_lock
	signal av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read                    : std_logic;                     -- av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> av_status_reg_0_avalon_slave_0_translator:uav_read
	signal av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata                : std_logic_vector(31 downto 0); -- av_status_reg_0_avalon_slave_0_translator:uav_readdata -> av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	signal av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid           : std_logic;                     -- av_status_reg_0_avalon_slave_0_translator:uav_readdatavalid -> av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess             : std_logic;                     -- av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> av_status_reg_0_avalon_slave_0_translator:uav_debugaccess
	signal av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable              : std_logic_vector(3 downto 0);  -- av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> av_status_reg_0_avalon_slave_0_translator:uav_byteenable
	signal av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket      : std_logic;                     -- av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid            : std_logic;                     -- av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket    : std_logic;                     -- av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data             : std_logic_vector(95 downto 0); -- av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready            : std_logic;                     -- av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket   : std_logic;                     -- av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid         : std_logic;                     -- av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket : std_logic;                     -- av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data          : std_logic_vector(95 downto 0); -- av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready         : std_logic;                     -- av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid       : std_logic;                     -- av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data        : std_logic_vector(33 downto 0); -- av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready       : std_logic;                     -- av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest             : std_logic;                     -- av_eth_config_0_avalon_slave_0_translator:uav_waitrequest -> av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount              : std_logic_vector(2 downto 0);  -- av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> av_eth_config_0_avalon_slave_0_translator:uav_burstcount
	signal av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata               : std_logic_vector(31 downto 0); -- av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> av_eth_config_0_avalon_slave_0_translator:uav_writedata
	signal av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address                 : std_logic_vector(19 downto 0); -- av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> av_eth_config_0_avalon_slave_0_translator:uav_address
	signal av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write                   : std_logic;                     -- av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> av_eth_config_0_avalon_slave_0_translator:uav_write
	signal av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock                    : std_logic;                     -- av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> av_eth_config_0_avalon_slave_0_translator:uav_lock
	signal av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read                    : std_logic;                     -- av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> av_eth_config_0_avalon_slave_0_translator:uav_read
	signal av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata                : std_logic_vector(31 downto 0); -- av_eth_config_0_avalon_slave_0_translator:uav_readdata -> av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	signal av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid           : std_logic;                     -- av_eth_config_0_avalon_slave_0_translator:uav_readdatavalid -> av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess             : std_logic;                     -- av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> av_eth_config_0_avalon_slave_0_translator:uav_debugaccess
	signal av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable              : std_logic_vector(3 downto 0);  -- av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> av_eth_config_0_avalon_slave_0_translator:uav_byteenable
	signal av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket      : std_logic;                     -- av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid            : std_logic;                     -- av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket    : std_logic;                     -- av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data             : std_logic_vector(95 downto 0); -- av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready            : std_logic;                     -- av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket   : std_logic;                     -- av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid         : std_logic;                     -- av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket : std_logic;                     -- av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data          : std_logic_vector(95 downto 0); -- av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready         : std_logic;                     -- av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid       : std_logic;                     -- av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data        : std_logic_vector(33 downto 0); -- av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready       : std_logic;                     -- av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest             : std_logic;                     -- av_config_reg_0_avalon_slave_0_translator:uav_waitrequest -> av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount              : std_logic_vector(2 downto 0);  -- av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> av_config_reg_0_avalon_slave_0_translator:uav_burstcount
	signal av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata               : std_logic_vector(31 downto 0); -- av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> av_config_reg_0_avalon_slave_0_translator:uav_writedata
	signal av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address                 : std_logic_vector(19 downto 0); -- av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> av_config_reg_0_avalon_slave_0_translator:uav_address
	signal av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write                   : std_logic;                     -- av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> av_config_reg_0_avalon_slave_0_translator:uav_write
	signal av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock                    : std_logic;                     -- av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> av_config_reg_0_avalon_slave_0_translator:uav_lock
	signal av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read                    : std_logic;                     -- av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> av_config_reg_0_avalon_slave_0_translator:uav_read
	signal av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata                : std_logic_vector(31 downto 0); -- av_config_reg_0_avalon_slave_0_translator:uav_readdata -> av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	signal av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid           : std_logic;                     -- av_config_reg_0_avalon_slave_0_translator:uav_readdatavalid -> av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess             : std_logic;                     -- av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> av_config_reg_0_avalon_slave_0_translator:uav_debugaccess
	signal av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable              : std_logic_vector(3 downto 0);  -- av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> av_config_reg_0_avalon_slave_0_translator:uav_byteenable
	signal av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket      : std_logic;                     -- av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid            : std_logic;                     -- av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket    : std_logic;                     -- av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data             : std_logic_vector(95 downto 0); -- av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready            : std_logic;                     -- av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket   : std_logic;                     -- av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid         : std_logic;                     -- av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket : std_logic;                     -- av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data          : std_logic_vector(95 downto 0); -- av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready         : std_logic;                     -- av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid       : std_logic;                     -- av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data        : std_logic_vector(33 downto 0); -- av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready       : std_logic;                     -- av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest             : std_logic;                     -- av_sendpacket_0_avalon_slave_0_translator:uav_waitrequest -> av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount              : std_logic_vector(2 downto 0);  -- av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> av_sendpacket_0_avalon_slave_0_translator:uav_burstcount
	signal av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata               : std_logic_vector(31 downto 0); -- av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> av_sendpacket_0_avalon_slave_0_translator:uav_writedata
	signal av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address                 : std_logic_vector(19 downto 0); -- av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> av_sendpacket_0_avalon_slave_0_translator:uav_address
	signal av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write                   : std_logic;                     -- av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> av_sendpacket_0_avalon_slave_0_translator:uav_write
	signal av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock                    : std_logic;                     -- av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> av_sendpacket_0_avalon_slave_0_translator:uav_lock
	signal av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read                    : std_logic;                     -- av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> av_sendpacket_0_avalon_slave_0_translator:uav_read
	signal av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata                : std_logic_vector(31 downto 0); -- av_sendpacket_0_avalon_slave_0_translator:uav_readdata -> av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	signal av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid           : std_logic;                     -- av_sendpacket_0_avalon_slave_0_translator:uav_readdatavalid -> av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess             : std_logic;                     -- av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> av_sendpacket_0_avalon_slave_0_translator:uav_debugaccess
	signal av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable              : std_logic_vector(3 downto 0);  -- av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> av_sendpacket_0_avalon_slave_0_translator:uav_byteenable
	signal av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket      : std_logic;                     -- av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid            : std_logic;                     -- av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket    : std_logic;                     -- av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data             : std_logic_vector(95 downto 0); -- av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready            : std_logic;                     -- av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket   : std_logic;                     -- av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid         : std_logic;                     -- av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket : std_logic;                     -- av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data          : std_logic_vector(95 downto 0); -- av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready         : std_logic;                     -- av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid       : std_logic;                     -- av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data        : std_logic_vector(33 downto 0); -- av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready       : std_logic;                     -- av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket           : std_logic;                     -- nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	signal nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid                 : std_logic;                     -- nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	signal nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket         : std_logic;                     -- nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	signal nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data                  : std_logic_vector(94 downto 0); -- nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	signal nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready                 : std_logic;                     -- addr_router:sink_ready -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	signal nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket                  : std_logic;                     -- nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	signal nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_valid                        : std_logic;                     -- nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	signal nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket                : std_logic;                     -- nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	signal nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_data                         : std_logic_vector(94 downto 0); -- nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	signal nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_ready                        : std_logic;                     -- addr_router_001:sink_ready -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_ready
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket             : std_logic;                     -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid                   : std_logic;                     -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket           : std_logic;                     -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data                    : std_logic_vector(94 downto 0); -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready                   : std_logic;                     -- id_router:sink_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                        : std_logic;                     -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_valid                              : std_logic;                     -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                      : std_logic;                     -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_data                               : std_logic_vector(94 downto 0); -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	signal onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_ready                              : std_logic;                     -- id_router_001:sink_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket              : std_logic;                     -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid                    : std_logic;                     -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket            : std_logic;                     -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data                     : std_logic_vector(94 downto 0); -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready                    : std_logic;                     -- id_router_002:sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket                 : std_logic;                     -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_valid                       : std_logic;                     -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket               : std_logic;                     -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_data                        : std_logic_vector(94 downto 0); -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_ready                       : std_logic;                     -- id_router_003:sink_ready -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                 : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid                                       : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                               : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data                                        : std_logic_vector(94 downto 0); -- timer_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready                                       : std_logic;                     -- id_router_004:sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal pio_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                   : std_logic;                     -- pio_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	signal pio_0_s1_translator_avalon_universal_slave_0_agent_rp_valid                                         : std_logic;                     -- pio_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	signal pio_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                 : std_logic;                     -- pio_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	signal pio_0_s1_translator_avalon_universal_slave_0_agent_rp_data                                          : std_logic_vector(94 downto 0); -- pio_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	signal pio_0_s1_translator_avalon_universal_slave_0_agent_rp_ready                                         : std_logic;                     -- id_router_005:sink_ready -> pio_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket             : std_logic;                     -- av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	signal av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid                   : std_logic;                     -- av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	signal av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket           : std_logic;                     -- av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	signal av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data                    : std_logic_vector(94 downto 0); -- av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	signal av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready                   : std_logic;                     -- id_router_006:sink_ready -> av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	signal av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket             : std_logic;                     -- av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	signal av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid                   : std_logic;                     -- av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	signal av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket           : std_logic;                     -- av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	signal av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data                    : std_logic_vector(94 downto 0); -- av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	signal av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready                   : std_logic;                     -- id_router_007:sink_ready -> av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	signal av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket             : std_logic;                     -- av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	signal av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid                   : std_logic;                     -- av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	signal av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket           : std_logic;                     -- av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	signal av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data                    : std_logic_vector(94 downto 0); -- av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	signal av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready                   : std_logic;                     -- id_router_008:sink_ready -> av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	signal av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket             : std_logic;                     -- av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	signal av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid                   : std_logic;                     -- av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	signal av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket           : std_logic;                     -- av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	signal av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data                    : std_logic_vector(94 downto 0); -- av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	signal av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready                   : std_logic;                     -- id_router_009:sink_ready -> av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	signal rst_controller_reset_out_reset                                                                      : std_logic;                     -- rst_controller:reset_out -> [addr_router:reset, addr_router_001:reset, av_config_reg_0_avalon_slave_0_translator:reset, av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, av_eth_config_0_avalon_slave_0_translator:reset, av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, av_sendpacket_0_avalon_slave_0_translator:reset, av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, av_status_reg_0_avalon_slave_0_translator:reset, av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, irq_mapper:reset, jtag_uart_0_avalon_jtag_slave_translator:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, nios2_qsys_0_data_master_translator:reset, nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:reset, nios2_qsys_0_instruction_master_translator:reset, nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:reset, nios2_qsys_0_jtag_debug_module_translator:reset, nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, onchip_memory2_0:reset, onchip_memory2_0_s1_translator:reset, onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:reset, onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_0_s1_translator:reset, pio_0_s1_translator_avalon_universal_slave_0_agent:reset, pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, rst_controller_reset_out_reset:in, sysid_qsys_0_control_slave_translator:reset, sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:reset, sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timer_0_s1_translator:reset, timer_0_s1_translator_avalon_universal_slave_0_agent:reset, timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	signal cmd_xbar_demux_src0_endofpacket                                                                     : std_logic;                     -- cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	signal cmd_xbar_demux_src0_valid                                                                           : std_logic;                     -- cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	signal cmd_xbar_demux_src0_startofpacket                                                                   : std_logic;                     -- cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	signal cmd_xbar_demux_src0_data                                                                            : std_logic_vector(94 downto 0); -- cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	signal cmd_xbar_demux_src0_channel                                                                         : std_logic_vector(9 downto 0);  -- cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	signal cmd_xbar_demux_src0_ready                                                                           : std_logic;                     -- cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	signal cmd_xbar_demux_src1_endofpacket                                                                     : std_logic;                     -- cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	signal cmd_xbar_demux_src1_valid                                                                           : std_logic;                     -- cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	signal cmd_xbar_demux_src1_startofpacket                                                                   : std_logic;                     -- cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	signal cmd_xbar_demux_src1_data                                                                            : std_logic_vector(94 downto 0); -- cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	signal cmd_xbar_demux_src1_channel                                                                         : std_logic_vector(9 downto 0);  -- cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	signal cmd_xbar_demux_src1_ready                                                                           : std_logic;                     -- cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	signal cmd_xbar_demux_001_src0_endofpacket                                                                 : std_logic;                     -- cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	signal cmd_xbar_demux_001_src0_valid                                                                       : std_logic;                     -- cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	signal cmd_xbar_demux_001_src0_startofpacket                                                               : std_logic;                     -- cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	signal cmd_xbar_demux_001_src0_data                                                                        : std_logic_vector(94 downto 0); -- cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	signal cmd_xbar_demux_001_src0_channel                                                                     : std_logic_vector(9 downto 0);  -- cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	signal cmd_xbar_demux_001_src0_ready                                                                       : std_logic;                     -- cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	signal cmd_xbar_demux_001_src1_endofpacket                                                                 : std_logic;                     -- cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	signal cmd_xbar_demux_001_src1_valid                                                                       : std_logic;                     -- cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	signal cmd_xbar_demux_001_src1_startofpacket                                                               : std_logic;                     -- cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	signal cmd_xbar_demux_001_src1_data                                                                        : std_logic_vector(94 downto 0); -- cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	signal cmd_xbar_demux_001_src1_channel                                                                     : std_logic_vector(9 downto 0);  -- cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	signal cmd_xbar_demux_001_src1_ready                                                                       : std_logic;                     -- cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	signal cmd_xbar_demux_001_src2_endofpacket                                                                 : std_logic;                     -- cmd_xbar_demux_001:src2_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src2_valid                                                                       : std_logic;                     -- cmd_xbar_demux_001:src2_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src2_startofpacket                                                               : std_logic;                     -- cmd_xbar_demux_001:src2_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src2_data                                                                        : std_logic_vector(94 downto 0); -- cmd_xbar_demux_001:src2_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src2_channel                                                                     : std_logic_vector(9 downto 0);  -- cmd_xbar_demux_001:src2_channel -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src3_endofpacket                                                                 : std_logic;                     -- cmd_xbar_demux_001:src3_endofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src3_valid                                                                       : std_logic;                     -- cmd_xbar_demux_001:src3_valid -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src3_startofpacket                                                               : std_logic;                     -- cmd_xbar_demux_001:src3_startofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src3_data                                                                        : std_logic_vector(94 downto 0); -- cmd_xbar_demux_001:src3_data -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src3_channel                                                                     : std_logic_vector(9 downto 0);  -- cmd_xbar_demux_001:src3_channel -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src4_endofpacket                                                                 : std_logic;                     -- cmd_xbar_demux_001:src4_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src4_valid                                                                       : std_logic;                     -- cmd_xbar_demux_001:src4_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src4_startofpacket                                                               : std_logic;                     -- cmd_xbar_demux_001:src4_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src4_data                                                                        : std_logic_vector(94 downto 0); -- cmd_xbar_demux_001:src4_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src4_channel                                                                     : std_logic_vector(9 downto 0);  -- cmd_xbar_demux_001:src4_channel -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src5_endofpacket                                                                 : std_logic;                     -- cmd_xbar_demux_001:src5_endofpacket -> pio_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src5_valid                                                                       : std_logic;                     -- cmd_xbar_demux_001:src5_valid -> pio_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src5_startofpacket                                                               : std_logic;                     -- cmd_xbar_demux_001:src5_startofpacket -> pio_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src5_data                                                                        : std_logic_vector(94 downto 0); -- cmd_xbar_demux_001:src5_data -> pio_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src5_channel                                                                     : std_logic_vector(9 downto 0);  -- cmd_xbar_demux_001:src5_channel -> pio_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src6_endofpacket                                                                 : std_logic;                     -- cmd_xbar_demux_001:src6_endofpacket -> av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src6_valid                                                                       : std_logic;                     -- cmd_xbar_demux_001:src6_valid -> av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src6_startofpacket                                                               : std_logic;                     -- cmd_xbar_demux_001:src6_startofpacket -> av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src6_data                                                                        : std_logic_vector(94 downto 0); -- cmd_xbar_demux_001:src6_data -> av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src6_channel                                                                     : std_logic_vector(9 downto 0);  -- cmd_xbar_demux_001:src6_channel -> av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src7_endofpacket                                                                 : std_logic;                     -- cmd_xbar_demux_001:src7_endofpacket -> av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src7_valid                                                                       : std_logic;                     -- cmd_xbar_demux_001:src7_valid -> av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src7_startofpacket                                                               : std_logic;                     -- cmd_xbar_demux_001:src7_startofpacket -> av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src7_data                                                                        : std_logic_vector(94 downto 0); -- cmd_xbar_demux_001:src7_data -> av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src7_channel                                                                     : std_logic_vector(9 downto 0);  -- cmd_xbar_demux_001:src7_channel -> av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src8_endofpacket                                                                 : std_logic;                     -- cmd_xbar_demux_001:src8_endofpacket -> av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src8_valid                                                                       : std_logic;                     -- cmd_xbar_demux_001:src8_valid -> av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src8_startofpacket                                                               : std_logic;                     -- cmd_xbar_demux_001:src8_startofpacket -> av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src8_data                                                                        : std_logic_vector(94 downto 0); -- cmd_xbar_demux_001:src8_data -> av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src8_channel                                                                     : std_logic_vector(9 downto 0);  -- cmd_xbar_demux_001:src8_channel -> av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src9_endofpacket                                                                 : std_logic;                     -- cmd_xbar_demux_001:src9_endofpacket -> av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src9_valid                                                                       : std_logic;                     -- cmd_xbar_demux_001:src9_valid -> av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src9_startofpacket                                                               : std_logic;                     -- cmd_xbar_demux_001:src9_startofpacket -> av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src9_data                                                                        : std_logic_vector(94 downto 0); -- cmd_xbar_demux_001:src9_data -> av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src9_channel                                                                     : std_logic_vector(9 downto 0);  -- cmd_xbar_demux_001:src9_channel -> av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	signal rsp_xbar_demux_src0_endofpacket                                                                     : std_logic;                     -- rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	signal rsp_xbar_demux_src0_valid                                                                           : std_logic;                     -- rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	signal rsp_xbar_demux_src0_startofpacket                                                                   : std_logic;                     -- rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	signal rsp_xbar_demux_src0_data                                                                            : std_logic_vector(94 downto 0); -- rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	signal rsp_xbar_demux_src0_channel                                                                         : std_logic_vector(9 downto 0);  -- rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	signal rsp_xbar_demux_src0_ready                                                                           : std_logic;                     -- rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	signal rsp_xbar_demux_src1_endofpacket                                                                     : std_logic;                     -- rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	signal rsp_xbar_demux_src1_valid                                                                           : std_logic;                     -- rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	signal rsp_xbar_demux_src1_startofpacket                                                                   : std_logic;                     -- rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	signal rsp_xbar_demux_src1_data                                                                            : std_logic_vector(94 downto 0); -- rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	signal rsp_xbar_demux_src1_channel                                                                         : std_logic_vector(9 downto 0);  -- rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	signal rsp_xbar_demux_src1_ready                                                                           : std_logic;                     -- rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	signal rsp_xbar_demux_001_src0_endofpacket                                                                 : std_logic;                     -- rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	signal rsp_xbar_demux_001_src0_valid                                                                       : std_logic;                     -- rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	signal rsp_xbar_demux_001_src0_startofpacket                                                               : std_logic;                     -- rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	signal rsp_xbar_demux_001_src0_data                                                                        : std_logic_vector(94 downto 0); -- rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	signal rsp_xbar_demux_001_src0_channel                                                                     : std_logic_vector(9 downto 0);  -- rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	signal rsp_xbar_demux_001_src0_ready                                                                       : std_logic;                     -- rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	signal rsp_xbar_demux_001_src1_endofpacket                                                                 : std_logic;                     -- rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	signal rsp_xbar_demux_001_src1_valid                                                                       : std_logic;                     -- rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	signal rsp_xbar_demux_001_src1_startofpacket                                                               : std_logic;                     -- rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	signal rsp_xbar_demux_001_src1_data                                                                        : std_logic_vector(94 downto 0); -- rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	signal rsp_xbar_demux_001_src1_channel                                                                     : std_logic_vector(9 downto 0);  -- rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	signal rsp_xbar_demux_001_src1_ready                                                                       : std_logic;                     -- rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	signal rsp_xbar_demux_002_src0_endofpacket                                                                 : std_logic;                     -- rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	signal rsp_xbar_demux_002_src0_valid                                                                       : std_logic;                     -- rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux_001:sink2_valid
	signal rsp_xbar_demux_002_src0_startofpacket                                                               : std_logic;                     -- rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	signal rsp_xbar_demux_002_src0_data                                                                        : std_logic_vector(94 downto 0); -- rsp_xbar_demux_002:src0_data -> rsp_xbar_mux_001:sink2_data
	signal rsp_xbar_demux_002_src0_channel                                                                     : std_logic_vector(9 downto 0);  -- rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux_001:sink2_channel
	signal rsp_xbar_demux_002_src0_ready                                                                       : std_logic;                     -- rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src0_ready
	signal rsp_xbar_demux_003_src0_endofpacket                                                                 : std_logic;                     -- rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	signal rsp_xbar_demux_003_src0_valid                                                                       : std_logic;                     -- rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux_001:sink3_valid
	signal rsp_xbar_demux_003_src0_startofpacket                                                               : std_logic;                     -- rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	signal rsp_xbar_demux_003_src0_data                                                                        : std_logic_vector(94 downto 0); -- rsp_xbar_demux_003:src0_data -> rsp_xbar_mux_001:sink3_data
	signal rsp_xbar_demux_003_src0_channel                                                                     : std_logic_vector(9 downto 0);  -- rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux_001:sink3_channel
	signal rsp_xbar_demux_003_src0_ready                                                                       : std_logic;                     -- rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src0_ready
	signal rsp_xbar_demux_004_src0_endofpacket                                                                 : std_logic;                     -- rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	signal rsp_xbar_demux_004_src0_valid                                                                       : std_logic;                     -- rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux_001:sink4_valid
	signal rsp_xbar_demux_004_src0_startofpacket                                                               : std_logic;                     -- rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	signal rsp_xbar_demux_004_src0_data                                                                        : std_logic_vector(94 downto 0); -- rsp_xbar_demux_004:src0_data -> rsp_xbar_mux_001:sink4_data
	signal rsp_xbar_demux_004_src0_channel                                                                     : std_logic_vector(9 downto 0);  -- rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux_001:sink4_channel
	signal rsp_xbar_demux_004_src0_ready                                                                       : std_logic;                     -- rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src0_ready
	signal rsp_xbar_demux_005_src0_endofpacket                                                                 : std_logic;                     -- rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	signal rsp_xbar_demux_005_src0_valid                                                                       : std_logic;                     -- rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux_001:sink5_valid
	signal rsp_xbar_demux_005_src0_startofpacket                                                               : std_logic;                     -- rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	signal rsp_xbar_demux_005_src0_data                                                                        : std_logic_vector(94 downto 0); -- rsp_xbar_demux_005:src0_data -> rsp_xbar_mux_001:sink5_data
	signal rsp_xbar_demux_005_src0_channel                                                                     : std_logic_vector(9 downto 0);  -- rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux_001:sink5_channel
	signal rsp_xbar_demux_005_src0_ready                                                                       : std_logic;                     -- rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_005:src0_ready
	signal rsp_xbar_demux_006_src0_endofpacket                                                                 : std_logic;                     -- rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	signal rsp_xbar_demux_006_src0_valid                                                                       : std_logic;                     -- rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux_001:sink6_valid
	signal rsp_xbar_demux_006_src0_startofpacket                                                               : std_logic;                     -- rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	signal rsp_xbar_demux_006_src0_data                                                                        : std_logic_vector(94 downto 0); -- rsp_xbar_demux_006:src0_data -> rsp_xbar_mux_001:sink6_data
	signal rsp_xbar_demux_006_src0_channel                                                                     : std_logic_vector(9 downto 0);  -- rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux_001:sink6_channel
	signal rsp_xbar_demux_006_src0_ready                                                                       : std_logic;                     -- rsp_xbar_mux_001:sink6_ready -> rsp_xbar_demux_006:src0_ready
	signal rsp_xbar_demux_007_src0_endofpacket                                                                 : std_logic;                     -- rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	signal rsp_xbar_demux_007_src0_valid                                                                       : std_logic;                     -- rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux_001:sink7_valid
	signal rsp_xbar_demux_007_src0_startofpacket                                                               : std_logic;                     -- rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	signal rsp_xbar_demux_007_src0_data                                                                        : std_logic_vector(94 downto 0); -- rsp_xbar_demux_007:src0_data -> rsp_xbar_mux_001:sink7_data
	signal rsp_xbar_demux_007_src0_channel                                                                     : std_logic_vector(9 downto 0);  -- rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux_001:sink7_channel
	signal rsp_xbar_demux_007_src0_ready                                                                       : std_logic;                     -- rsp_xbar_mux_001:sink7_ready -> rsp_xbar_demux_007:src0_ready
	signal rsp_xbar_demux_008_src0_endofpacket                                                                 : std_logic;                     -- rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux_001:sink8_endofpacket
	signal rsp_xbar_demux_008_src0_valid                                                                       : std_logic;                     -- rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux_001:sink8_valid
	signal rsp_xbar_demux_008_src0_startofpacket                                                               : std_logic;                     -- rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux_001:sink8_startofpacket
	signal rsp_xbar_demux_008_src0_data                                                                        : std_logic_vector(94 downto 0); -- rsp_xbar_demux_008:src0_data -> rsp_xbar_mux_001:sink8_data
	signal rsp_xbar_demux_008_src0_channel                                                                     : std_logic_vector(9 downto 0);  -- rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux_001:sink8_channel
	signal rsp_xbar_demux_008_src0_ready                                                                       : std_logic;                     -- rsp_xbar_mux_001:sink8_ready -> rsp_xbar_demux_008:src0_ready
	signal rsp_xbar_demux_009_src0_endofpacket                                                                 : std_logic;                     -- rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux_001:sink9_endofpacket
	signal rsp_xbar_demux_009_src0_valid                                                                       : std_logic;                     -- rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux_001:sink9_valid
	signal rsp_xbar_demux_009_src0_startofpacket                                                               : std_logic;                     -- rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux_001:sink9_startofpacket
	signal rsp_xbar_demux_009_src0_data                                                                        : std_logic_vector(94 downto 0); -- rsp_xbar_demux_009:src0_data -> rsp_xbar_mux_001:sink9_data
	signal rsp_xbar_demux_009_src0_channel                                                                     : std_logic_vector(9 downto 0);  -- rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux_001:sink9_channel
	signal rsp_xbar_demux_009_src0_ready                                                                       : std_logic;                     -- rsp_xbar_mux_001:sink9_ready -> rsp_xbar_demux_009:src0_ready
	signal addr_router_src_endofpacket                                                                         : std_logic;                     -- addr_router:src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	signal addr_router_src_valid                                                                               : std_logic;                     -- addr_router:src_valid -> cmd_xbar_demux:sink_valid
	signal addr_router_src_startofpacket                                                                       : std_logic;                     -- addr_router:src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	signal addr_router_src_data                                                                                : std_logic_vector(94 downto 0); -- addr_router:src_data -> cmd_xbar_demux:sink_data
	signal addr_router_src_channel                                                                             : std_logic_vector(9 downto 0);  -- addr_router:src_channel -> cmd_xbar_demux:sink_channel
	signal addr_router_src_ready                                                                               : std_logic;                     -- cmd_xbar_demux:sink_ready -> addr_router:src_ready
	signal rsp_xbar_mux_src_endofpacket                                                                        : std_logic;                     -- rsp_xbar_mux:src_endofpacket -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal rsp_xbar_mux_src_valid                                                                              : std_logic;                     -- rsp_xbar_mux:src_valid -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	signal rsp_xbar_mux_src_startofpacket                                                                      : std_logic;                     -- rsp_xbar_mux:src_startofpacket -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal rsp_xbar_mux_src_data                                                                               : std_logic_vector(94 downto 0); -- rsp_xbar_mux:src_data -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	signal rsp_xbar_mux_src_channel                                                                            : std_logic_vector(9 downto 0);  -- rsp_xbar_mux:src_channel -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	signal rsp_xbar_mux_src_ready                                                                              : std_logic;                     -- nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux:src_ready
	signal addr_router_001_src_endofpacket                                                                     : std_logic;                     -- addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	signal addr_router_001_src_valid                                                                           : std_logic;                     -- addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	signal addr_router_001_src_startofpacket                                                                   : std_logic;                     -- addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	signal addr_router_001_src_data                                                                            : std_logic_vector(94 downto 0); -- addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	signal addr_router_001_src_channel                                                                         : std_logic_vector(9 downto 0);  -- addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	signal addr_router_001_src_ready                                                                           : std_logic;                     -- cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	signal rsp_xbar_mux_001_src_endofpacket                                                                    : std_logic;                     -- rsp_xbar_mux_001:src_endofpacket -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal rsp_xbar_mux_001_src_valid                                                                          : std_logic;                     -- rsp_xbar_mux_001:src_valid -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_valid
	signal rsp_xbar_mux_001_src_startofpacket                                                                  : std_logic;                     -- rsp_xbar_mux_001:src_startofpacket -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal rsp_xbar_mux_001_src_data                                                                           : std_logic_vector(94 downto 0); -- rsp_xbar_mux_001:src_data -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_data
	signal rsp_xbar_mux_001_src_channel                                                                        : std_logic_vector(9 downto 0);  -- rsp_xbar_mux_001:src_channel -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_channel
	signal rsp_xbar_mux_001_src_ready                                                                          : std_logic;                     -- nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_001:src_ready
	signal cmd_xbar_mux_src_endofpacket                                                                        : std_logic;                     -- cmd_xbar_mux:src_endofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_src_valid                                                                              : std_logic;                     -- cmd_xbar_mux:src_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_src_startofpacket                                                                      : std_logic;                     -- cmd_xbar_mux:src_startofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_src_data                                                                               : std_logic_vector(94 downto 0); -- cmd_xbar_mux:src_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_src_channel                                                                            : std_logic_vector(9 downto 0);  -- cmd_xbar_mux:src_channel -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_src_ready                                                                              : std_logic;                     -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	signal id_router_src_endofpacket                                                                           : std_logic;                     -- id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	signal id_router_src_valid                                                                                 : std_logic;                     -- id_router:src_valid -> rsp_xbar_demux:sink_valid
	signal id_router_src_startofpacket                                                                         : std_logic;                     -- id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	signal id_router_src_data                                                                                  : std_logic_vector(94 downto 0); -- id_router:src_data -> rsp_xbar_demux:sink_data
	signal id_router_src_channel                                                                               : std_logic_vector(9 downto 0);  -- id_router:src_channel -> rsp_xbar_demux:sink_channel
	signal id_router_src_ready                                                                                 : std_logic;                     -- rsp_xbar_demux:sink_ready -> id_router:src_ready
	signal cmd_xbar_mux_001_src_endofpacket                                                                    : std_logic;                     -- cmd_xbar_mux_001:src_endofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_001_src_valid                                                                          : std_logic;                     -- cmd_xbar_mux_001:src_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_001_src_startofpacket                                                                  : std_logic;                     -- cmd_xbar_mux_001:src_startofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_001_src_data                                                                           : std_logic_vector(94 downto 0); -- cmd_xbar_mux_001:src_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_001_src_channel                                                                        : std_logic_vector(9 downto 0);  -- cmd_xbar_mux_001:src_channel -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_001_src_ready                                                                          : std_logic;                     -- onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_001:src_ready
	signal id_router_001_src_endofpacket                                                                       : std_logic;                     -- id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	signal id_router_001_src_valid                                                                             : std_logic;                     -- id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	signal id_router_001_src_startofpacket                                                                     : std_logic;                     -- id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	signal id_router_001_src_data                                                                              : std_logic_vector(94 downto 0); -- id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	signal id_router_001_src_channel                                                                           : std_logic_vector(9 downto 0);  -- id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	signal id_router_001_src_ready                                                                             : std_logic;                     -- rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	signal cmd_xbar_demux_001_src2_ready                                                                       : std_logic;                     -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src2_ready
	signal id_router_002_src_endofpacket                                                                       : std_logic;                     -- id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	signal id_router_002_src_valid                                                                             : std_logic;                     -- id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	signal id_router_002_src_startofpacket                                                                     : std_logic;                     -- id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	signal id_router_002_src_data                                                                              : std_logic_vector(94 downto 0); -- id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	signal id_router_002_src_channel                                                                           : std_logic_vector(9 downto 0);  -- id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	signal id_router_002_src_ready                                                                             : std_logic;                     -- rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	signal cmd_xbar_demux_001_src3_ready                                                                       : std_logic;                     -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src3_ready
	signal id_router_003_src_endofpacket                                                                       : std_logic;                     -- id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	signal id_router_003_src_valid                                                                             : std_logic;                     -- id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	signal id_router_003_src_startofpacket                                                                     : std_logic;                     -- id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	signal id_router_003_src_data                                                                              : std_logic_vector(94 downto 0); -- id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	signal id_router_003_src_channel                                                                           : std_logic_vector(9 downto 0);  -- id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	signal id_router_003_src_ready                                                                             : std_logic;                     -- rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	signal cmd_xbar_demux_001_src4_ready                                                                       : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src4_ready
	signal id_router_004_src_endofpacket                                                                       : std_logic;                     -- id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	signal id_router_004_src_valid                                                                             : std_logic;                     -- id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	signal id_router_004_src_startofpacket                                                                     : std_logic;                     -- id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	signal id_router_004_src_data                                                                              : std_logic_vector(94 downto 0); -- id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	signal id_router_004_src_channel                                                                           : std_logic_vector(9 downto 0);  -- id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	signal id_router_004_src_ready                                                                             : std_logic;                     -- rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	signal cmd_xbar_demux_001_src5_ready                                                                       : std_logic;                     -- pio_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src5_ready
	signal id_router_005_src_endofpacket                                                                       : std_logic;                     -- id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	signal id_router_005_src_valid                                                                             : std_logic;                     -- id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	signal id_router_005_src_startofpacket                                                                     : std_logic;                     -- id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	signal id_router_005_src_data                                                                              : std_logic_vector(94 downto 0); -- id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	signal id_router_005_src_channel                                                                           : std_logic_vector(9 downto 0);  -- id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	signal id_router_005_src_ready                                                                             : std_logic;                     -- rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	signal cmd_xbar_demux_001_src6_ready                                                                       : std_logic;                     -- av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src6_ready
	signal id_router_006_src_endofpacket                                                                       : std_logic;                     -- id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	signal id_router_006_src_valid                                                                             : std_logic;                     -- id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	signal id_router_006_src_startofpacket                                                                     : std_logic;                     -- id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	signal id_router_006_src_data                                                                              : std_logic_vector(94 downto 0); -- id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	signal id_router_006_src_channel                                                                           : std_logic_vector(9 downto 0);  -- id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	signal id_router_006_src_ready                                                                             : std_logic;                     -- rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	signal cmd_xbar_demux_001_src7_ready                                                                       : std_logic;                     -- av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src7_ready
	signal id_router_007_src_endofpacket                                                                       : std_logic;                     -- id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	signal id_router_007_src_valid                                                                             : std_logic;                     -- id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	signal id_router_007_src_startofpacket                                                                     : std_logic;                     -- id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	signal id_router_007_src_data                                                                              : std_logic_vector(94 downto 0); -- id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	signal id_router_007_src_channel                                                                           : std_logic_vector(9 downto 0);  -- id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	signal id_router_007_src_ready                                                                             : std_logic;                     -- rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	signal cmd_xbar_demux_001_src8_ready                                                                       : std_logic;                     -- av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src8_ready
	signal id_router_008_src_endofpacket                                                                       : std_logic;                     -- id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	signal id_router_008_src_valid                                                                             : std_logic;                     -- id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	signal id_router_008_src_startofpacket                                                                     : std_logic;                     -- id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	signal id_router_008_src_data                                                                              : std_logic_vector(94 downto 0); -- id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	signal id_router_008_src_channel                                                                           : std_logic_vector(9 downto 0);  -- id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	signal id_router_008_src_ready                                                                             : std_logic;                     -- rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	signal cmd_xbar_demux_001_src9_ready                                                                       : std_logic;                     -- av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src9_ready
	signal id_router_009_src_endofpacket                                                                       : std_logic;                     -- id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	signal id_router_009_src_valid                                                                             : std_logic;                     -- id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	signal id_router_009_src_startofpacket                                                                     : std_logic;                     -- id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	signal id_router_009_src_data                                                                              : std_logic_vector(94 downto 0); -- id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	signal id_router_009_src_channel                                                                           : std_logic_vector(9 downto 0);  -- id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	signal id_router_009_src_ready                                                                             : std_logic;                     -- rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	signal irq_mapper_receiver0_irq                                                                            : std_logic;                     -- timer_0:irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                                                            : std_logic;                     -- jtag_uart_0:av_irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                                                            : std_logic;                     -- av_config_reg_0:av_irq -> irq_mapper:receiver2_irq
	signal nios2_qsys_0_d_irq_irq                                                                              : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2_qsys_0:d_irq
	signal reset_reset_n_ports_inv                                                                             : std_logic;                     -- reset_reset_n:inv -> rst_controller:reset_in0
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write_ports_inv                        : std_logic;                     -- jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write:inv -> jtag_uart_0:av_write_n
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read_ports_inv                         : std_logic;                     -- jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read:inv -> jtag_uart_0:av_read_n
	signal timer_0_s1_translator_avalon_anti_slave_0_write_ports_inv                                           : std_logic;                     -- timer_0_s1_translator_avalon_anti_slave_0_write:inv -> timer_0:write_n
	signal pio_0_s1_translator_avalon_anti_slave_0_write_ports_inv                                             : std_logic;                     -- pio_0_s1_translator_avalon_anti_slave_0_write:inv -> pio_0:write_n
	signal rst_controller_reset_out_reset_ports_inv                                                            : std_logic;                     -- rst_controller_reset_out_reset:inv -> [av_config_reg_0:reset_n, av_eth_config_0:reset_n, av_sendpacket_0:reset_n, av_status_reg_0:reset_n, jtag_uart_0:rst_n, nios2_qsys_0:reset_n, pio_0:reset_n, sysid_qsys_0:reset_n, timer_0:reset_n]

begin

	onchip_memory2_0 : component nios_system_onchip_memory2_0
		port map (
			clk        => clk_clk,                                                       --   clk1.clk
			address    => onchip_memory2_0_s1_translator_avalon_anti_slave_0_address,    --     s1.address
			clken      => onchip_memory2_0_s1_translator_avalon_anti_slave_0_clken,      --       .clken
			chipselect => onchip_memory2_0_s1_translator_avalon_anti_slave_0_chipselect, --       .chipselect
			write      => onchip_memory2_0_s1_translator_avalon_anti_slave_0_write,      --       .write
			readdata   => onchip_memory2_0_s1_translator_avalon_anti_slave_0_readdata,   --       .readdata
			writedata  => onchip_memory2_0_s1_translator_avalon_anti_slave_0_writedata,  --       .writedata
			byteenable => onchip_memory2_0_s1_translator_avalon_anti_slave_0_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset                                 -- reset1.reset
		);

	nios2_qsys_0 : component nios_system_nios2_qsys_0
		port map (
			clk                                   => clk_clk,                                                                   --                       clk.clk
			reset_n                               => rst_controller_reset_out_reset_ports_inv,                                  --                   reset_n.reset_n
			d_address                             => nios2_qsys_0_data_master_address,                                          --               data_master.address
			d_byteenable                          => nios2_qsys_0_data_master_byteenable,                                       --                          .byteenable
			d_read                                => nios2_qsys_0_data_master_read,                                             --                          .read
			d_readdata                            => nios2_qsys_0_data_master_readdata,                                         --                          .readdata
			d_waitrequest                         => nios2_qsys_0_data_master_waitrequest,                                      --                          .waitrequest
			d_write                               => nios2_qsys_0_data_master_write,                                            --                          .write
			d_writedata                           => nios2_qsys_0_data_master_writedata,                                        --                          .writedata
			jtag_debug_module_debugaccess_to_roms => nios2_qsys_0_data_master_debugaccess,                                      --                          .debugaccess
			i_address                             => nios2_qsys_0_instruction_master_address,                                   --        instruction_master.address
			i_read                                => nios2_qsys_0_instruction_master_read,                                      --                          .read
			i_readdata                            => nios2_qsys_0_instruction_master_readdata,                                  --                          .readdata
			i_waitrequest                         => nios2_qsys_0_instruction_master_waitrequest,                               --                          .waitrequest
			d_irq                                 => nios2_qsys_0_d_irq_irq,                                                    --                     d_irq.irq
			jtag_debug_module_resetrequest        => open,                                                                      --   jtag_debug_module_reset.reset
			jtag_debug_module_address             => nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_address,     --         jtag_debug_module.address
			jtag_debug_module_byteenable          => nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable,  --                          .byteenable
			jtag_debug_module_debugaccess         => nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess, --                          .debugaccess
			jtag_debug_module_read                => nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_read,        --                          .read
			jtag_debug_module_readdata            => nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata,    --                          .readdata
			jtag_debug_module_waitrequest         => nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest, --                          .waitrequest
			jtag_debug_module_write               => nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_write,       --                          .write
			jtag_debug_module_writedata           => nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata,   --                          .writedata
			no_ci_readra                          => open                                                                       -- custom_instruction_master.readra
		);

	jtag_uart_0 : component nios_system_jtag_uart_0
		port map (
			clk            => clk_clk,                                                                      --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                                     --             reset.reset_n
			av_chipselect  => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address(0),      --                  .address
			av_read_n      => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read_ports_inv,  --                  .read_n
			av_readdata    => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata,        --                  .readdata
			av_write_n     => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write_ports_inv, --                  .write_n
			av_writedata   => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata,       --                  .writedata
			av_waitrequest => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver1_irq                                                      --               irq.irq
		);

	sysid_qsys_0 : component nios_system_sysid_qsys_0
		port map (
			clock    => clk_clk,                                                              --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,                             --         reset.reset_n
			readdata => sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_readdata,   -- control_slave.readdata
			address  => sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_address(0)  --              .address
		);

	timer_0 : component nios_system_timer_0
		port map (
			clk        => clk_clk,                                                   --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                  -- reset.reset_n
			address    => timer_0_s1_translator_avalon_anti_slave_0_address,         --    s1.address
			writedata  => timer_0_s1_translator_avalon_anti_slave_0_writedata,       --      .writedata
			readdata   => timer_0_s1_translator_avalon_anti_slave_0_readdata,        --      .readdata
			chipselect => timer_0_s1_translator_avalon_anti_slave_0_chipselect,      --      .chipselect
			write_n    => timer_0_s1_translator_avalon_anti_slave_0_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver0_irq                                   --   irq.irq
		);

	pio_0 : component nios_system_pio_0
		port map (
			clk        => clk_clk,                                                 --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                --               reset.reset_n
			address    => pio_0_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => pio_0_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => pio_0_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => pio_0_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => pio_0_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => pio_0_external_connection_export                         -- external_connection.export
		);

	av_status_reg_0 : component av_status_reg
		port map (
			clk           => clk_clk,                                                                 --          clock.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,                                --          reset.reset_n
			address       => av_status_reg_0_avalon_slave_0_translator_avalon_anti_slave_0_address,   -- avalon_slave_0.address
			write         => av_status_reg_0_avalon_slave_0_translator_avalon_anti_slave_0_write,     --               .write
			read          => av_status_reg_0_avalon_slave_0_translator_avalon_anti_slave_0_read,      --               .read
			writedata     => av_status_reg_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata, --               .writedata
			readdata      => av_status_reg_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata,  --               .readdata
			udp_send      => av_status_reg_0_conduit_end_udp_send,                                    --    conduit_end.export
			status_reg0_o => av_status_reg_0_conduit_end_status_reg0_o,                               --               .export
			status_reg1_o => av_status_reg_0_conduit_end_status_reg1_o,                               --               .export
			status_reg2_o => av_status_reg_0_conduit_end_status_reg2_o,                               --               .export
			status_reg3_o => av_status_reg_0_conduit_end_status_reg3_o,                               --               .export
			status_reg4_o => av_status_reg_0_conduit_end_status_reg4_o,                               --               .export
			status_reg5_o => av_status_reg_0_conduit_end_status_reg5_o,                               --               .export
			status_reg7_o => av_status_reg_0_conduit_end_status_reg7_o,                               --               .export
			status_reg6_o => av_status_reg_0_conduit_end_status_reg6_o                                --               .export
		);

	av_eth_config_0 : component av_eth_config
		port map (
			clk              => clk_clk,                                                                 --          clock.clk
			reset_n          => rst_controller_reset_out_reset_ports_inv,                                --          reset.reset_n
			write            => av_eth_config_0_avalon_slave_0_translator_avalon_anti_slave_0_write,     -- avalon_slave_0.write
			read             => av_eth_config_0_avalon_slave_0_translator_avalon_anti_slave_0_read,      --               .read
			writedata        => av_eth_config_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata, --               .writedata
			address          => av_eth_config_0_avalon_slave_0_translator_avalon_anti_slave_0_address,   --               .address
			readdata         => av_eth_config_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata,  --               .readdata
			local_port_o     => av_eth_config_0_conduit_end_local_port_o,                                --    conduit_end.export
			remote_port_o    => av_eth_config_0_conduit_end_remote_port_o,                               --               .export
			local_IP_o       => av_eth_config_0_conduit_end_local_IP_o,                                  --               .export
			remote_IP_o      => av_eth_config_0_conduit_end_remote_IP_o,                                 --               .export
			local_MAC_LSB_o  => av_eth_config_0_conduit_end_local_MAC_LSB_o,                             --               .export
			local_MAC_MSB_o  => av_eth_config_0_conduit_end_local_MAC_MSB_o,                             --               .export
			remote_MAC_LSB_o => av_eth_config_0_conduit_end_remote_MAC_LSB_o,                            --               .export
			checksum_o       => av_eth_config_0_conduit_end_checksum_o,                                  --               .export
			remote_MAC_MSB_o => av_eth_config_0_conduit_end_remote_MAC_MSB_o                             --               .export
		);

	av_config_reg_0 : component av_config_reg
		port map (
			clk            => clk_clk,                                                                 --            clock.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,                                --            reset.reset_n
			address        => av_config_reg_0_avalon_slave_0_translator_avalon_anti_slave_0_address,   --   avalon_slave_0.address
			write          => av_config_reg_0_avalon_slave_0_translator_avalon_anti_slave_0_write,     --                 .write
			read           => av_config_reg_0_avalon_slave_0_translator_avalon_anti_slave_0_read,      --                 .read
			writedata      => av_config_reg_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata, --                 .writedata
			readdata       => av_config_reg_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata,  --                 .readdata
			reg_0          => av_config_reg_0_conduit_end_reg_0,                                       --      conduit_end.export
			reg_1          => av_config_reg_0_conduit_end_reg_1,                                       --                 .export
			reg_2          => av_config_reg_0_conduit_end_reg_2,                                       --                 .export
			reg_3          => av_config_reg_0_conduit_end_reg_3,                                       --                 .export
			reg_4          => av_config_reg_0_conduit_end_reg_4,                                       --                 .export
			reg_5          => av_config_reg_0_conduit_end_reg_5,                                       --                 .export
			reg_6          => av_config_reg_0_conduit_end_reg_6,                                       --                 .export
			reg_7          => av_config_reg_0_conduit_end_reg_7,                                       --                 .export
			udp_data_valid => av_config_reg_0_conduit_end_udp_data_valid,                              --                 .export
			av_irq         => irq_mapper_receiver2_irq                                                 -- interrupt_sender.irq
		);

	av_sendpacket_0 : component av_sendpacket
		port map (
			clk              => clk_clk,                                                                 --          clock.clk
			reset_n          => rst_controller_reset_out_reset_ports_inv,                                --          reset.reset_n
			address          => av_sendpacket_0_avalon_slave_0_translator_avalon_anti_slave_0_address,   -- avalon_slave_0.address
			write            => av_sendpacket_0_avalon_slave_0_translator_avalon_anti_slave_0_write,     --               .write
			read             => av_sendpacket_0_avalon_slave_0_translator_avalon_anti_slave_0_read,      --               .read
			writedata        => av_sendpacket_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata, --               .writedata
			readdata         => av_sendpacket_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata,  --               .readdata
			checksum_o       => av_sendpacket_0_conduit_end_checksum_o,                                  --    conduit_end.export
			local_port_o     => av_sendpacket_0_conduit_end_local_port_o,                                --               .export
			remote_port_o    => av_sendpacket_0_conduit_end_remote_port_o,                               --               .export
			remote_MAC_MSB_o => av_sendpacket_0_conduit_end_remote_MAC_MSB_o,                            --               .export
			remote_MAC_LSB_o => av_sendpacket_0_conduit_end_remote_MAC_LSB_o,                            --               .export
			udp_sendpacket   => av_sendpacket_0_conduit_end_udp_sendpacket,                              --               .export
			length_o         => av_sendpacket_0_conduit_end_length_o,                                    --               .export
			remote_IP_o      => av_sendpacket_0_conduit_end_remote_IP_o                                  --               .export
		);

	nios2_qsys_0_instruction_master_translator : component nios_system_nios2_qsys_0_instruction_master_translator
		generic map (
			AV_ADDRESS_W                => 20,
			AV_DATA_W                   => 32,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 4,
			UAV_ADDRESS_W               => 20,
			UAV_BURSTCOUNT_W            => 3,
			USE_READ                    => 1,
			USE_WRITE                   => 0,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 0,
			USE_READDATAVALID           => 0,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 4,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 1,
			AV_REGISTERINCOMINGSIGNALS  => 0
		)
		port map (
			clk                      => clk_clk,                                                                            --                       clk.clk
			reset                    => rst_controller_reset_out_reset,                                                     --                     reset.reset
			uav_address              => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => nios2_qsys_0_instruction_master_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => nios2_qsys_0_instruction_master_waitrequest,                                        --                          .waitrequest
			av_read                  => nios2_qsys_0_instruction_master_read,                                               --                          .read
			av_readdata              => nios2_qsys_0_instruction_master_readdata,                                           --                          .readdata
			av_burstcount            => "1",                                                                                --               (terminated)
			av_byteenable            => "1111",                                                                             --               (terminated)
			av_beginbursttransfer    => '0',                                                                                --               (terminated)
			av_begintransfer         => '0',                                                                                --               (terminated)
			av_chipselect            => '0',                                                                                --               (terminated)
			av_readdatavalid         => open,                                                                               --               (terminated)
			av_write                 => '0',                                                                                --               (terminated)
			av_writedata             => "00000000000000000000000000000000",                                                 --               (terminated)
			av_lock                  => '0',                                                                                --               (terminated)
			av_debugaccess           => '0',                                                                                --               (terminated)
			uav_clken                => open,                                                                               --               (terminated)
			av_clken                 => '1',                                                                                --               (terminated)
			uav_response             => "00",                                                                               --               (terminated)
			av_response              => open,                                                                               --               (terminated)
			uav_writeresponserequest => open,                                                                               --               (terminated)
			uav_writeresponsevalid   => '0',                                                                                --               (terminated)
			av_writeresponserequest  => '0',                                                                                --               (terminated)
			av_writeresponsevalid    => open                                                                                --               (terminated)
		);

	nios2_qsys_0_data_master_translator : component nios_system_nios2_qsys_0_data_master_translator
		generic map (
			AV_ADDRESS_W                => 20,
			AV_DATA_W                   => 32,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 4,
			UAV_ADDRESS_W               => 20,
			UAV_BURSTCOUNT_W            => 3,
			USE_READ                    => 1,
			USE_WRITE                   => 1,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 0,
			USE_READDATAVALID           => 0,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 4,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 0,
			AV_REGISTERINCOMINGSIGNALS  => 1
		)
		port map (
			clk                      => clk_clk,                                                                     --                       clk.clk
			reset                    => rst_controller_reset_out_reset,                                              --                     reset.reset
			uav_address              => nios2_qsys_0_data_master_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => nios2_qsys_0_data_master_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => nios2_qsys_0_data_master_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => nios2_qsys_0_data_master_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => nios2_qsys_0_data_master_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => nios2_qsys_0_data_master_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => nios2_qsys_0_data_master_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => nios2_qsys_0_data_master_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => nios2_qsys_0_data_master_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => nios2_qsys_0_data_master_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => nios2_qsys_0_data_master_waitrequest,                                        --                          .waitrequest
			av_byteenable            => nios2_qsys_0_data_master_byteenable,                                         --                          .byteenable
			av_read                  => nios2_qsys_0_data_master_read,                                               --                          .read
			av_readdata              => nios2_qsys_0_data_master_readdata,                                           --                          .readdata
			av_write                 => nios2_qsys_0_data_master_write,                                              --                          .write
			av_writedata             => nios2_qsys_0_data_master_writedata,                                          --                          .writedata
			av_debugaccess           => nios2_qsys_0_data_master_debugaccess,                                        --                          .debugaccess
			av_burstcount            => "1",                                                                         --               (terminated)
			av_beginbursttransfer    => '0',                                                                         --               (terminated)
			av_begintransfer         => '0',                                                                         --               (terminated)
			av_chipselect            => '0',                                                                         --               (terminated)
			av_readdatavalid         => open,                                                                        --               (terminated)
			av_lock                  => '0',                                                                         --               (terminated)
			uav_clken                => open,                                                                        --               (terminated)
			av_clken                 => '1',                                                                         --               (terminated)
			uav_response             => "00",                                                                        --               (terminated)
			av_response              => open,                                                                        --               (terminated)
			uav_writeresponserequest => open,                                                                        --               (terminated)
			uav_writeresponsevalid   => '0',                                                                         --               (terminated)
			av_writeresponserequest  => '0',                                                                         --               (terminated)
			av_writeresponsevalid    => open                                                                         --               (terminated)
		);

	nios2_qsys_0_jtag_debug_module_translator : component nios_system_nios2_qsys_0_jtag_debug_module_translator
		generic map (
			AV_ADDRESS_W                   => 9,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 20,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                                                   --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                            --                    reset.reset
			uav_address              => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_waitrequest           => nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_debugaccess           => nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess,                 --                         .debugaccess
			av_begintransfer         => open,                                                                                      --              (terminated)
			av_beginbursttransfer    => open,                                                                                      --              (terminated)
			av_burstcount            => open,                                                                                      --              (terminated)
			av_readdatavalid         => '0',                                                                                       --              (terminated)
			av_writebyteenable       => open,                                                                                      --              (terminated)
			av_lock                  => open,                                                                                      --              (terminated)
			av_chipselect            => open,                                                                                      --              (terminated)
			av_clken                 => open,                                                                                      --              (terminated)
			uav_clken                => '0',                                                                                       --              (terminated)
			av_outputenable          => open,                                                                                      --              (terminated)
			uav_response             => open,                                                                                      --              (terminated)
			av_response              => "00",                                                                                      --              (terminated)
			uav_writeresponserequest => '0',                                                                                       --              (terminated)
			uav_writeresponsevalid   => open,                                                                                      --              (terminated)
			av_writeresponserequest  => open,                                                                                      --              (terminated)
			av_writeresponsevalid    => '0'                                                                                        --              (terminated)
		);

	onchip_memory2_0_s1_translator : component nios_system_onchip_memory2_0_s1_translator
		generic map (
			AV_ADDRESS_W                   => 16,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 20,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 1,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 0,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                                        --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                 --                    reset.reset
			uav_address              => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => onchip_memory2_0_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => onchip_memory2_0_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => onchip_memory2_0_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => onchip_memory2_0_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => onchip_memory2_0_s1_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_chipselect            => onchip_memory2_0_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_clken                 => onchip_memory2_0_s1_translator_avalon_anti_slave_0_clken,                       --                         .clken
			av_read                  => open,                                                                           --              (terminated)
			av_begintransfer         => open,                                                                           --              (terminated)
			av_beginbursttransfer    => open,                                                                           --              (terminated)
			av_burstcount            => open,                                                                           --              (terminated)
			av_readdatavalid         => '0',                                                                            --              (terminated)
			av_waitrequest           => '0',                                                                            --              (terminated)
			av_writebyteenable       => open,                                                                           --              (terminated)
			av_lock                  => open,                                                                           --              (terminated)
			uav_clken                => '0',                                                                            --              (terminated)
			av_debugaccess           => open,                                                                           --              (terminated)
			av_outputenable          => open,                                                                           --              (terminated)
			uav_response             => open,                                                                           --              (terminated)
			av_response              => "00",                                                                           --              (terminated)
			uav_writeresponserequest => '0',                                                                            --              (terminated)
			uav_writeresponsevalid   => open,                                                                           --              (terminated)
			av_writeresponserequest  => open,                                                                           --              (terminated)
			av_writeresponsevalid    => '0'                                                                             --              (terminated)
		);

	jtag_uart_0_avalon_jtag_slave_translator : component nios_system_jtag_uart_0_avalon_jtag_slave_translator
		generic map (
			AV_ADDRESS_W                   => 1,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 20,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                                                  --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                           --                    reset.reset
			uav_address              => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_waitrequest           => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_chipselect            => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_begintransfer         => open,                                                                                     --              (terminated)
			av_beginbursttransfer    => open,                                                                                     --              (terminated)
			av_burstcount            => open,                                                                                     --              (terminated)
			av_byteenable            => open,                                                                                     --              (terminated)
			av_readdatavalid         => '0',                                                                                      --              (terminated)
			av_writebyteenable       => open,                                                                                     --              (terminated)
			av_lock                  => open,                                                                                     --              (terminated)
			av_clken                 => open,                                                                                     --              (terminated)
			uav_clken                => '0',                                                                                      --              (terminated)
			av_debugaccess           => open,                                                                                     --              (terminated)
			av_outputenable          => open,                                                                                     --              (terminated)
			uav_response             => open,                                                                                     --              (terminated)
			av_response              => "00",                                                                                     --              (terminated)
			uav_writeresponserequest => '0',                                                                                      --              (terminated)
			uav_writeresponsevalid   => open,                                                                                     --              (terminated)
			av_writeresponserequest  => open,                                                                                     --              (terminated)
			av_writeresponsevalid    => '0'                                                                                       --              (terminated)
		);

	sysid_qsys_0_control_slave_translator : component nios_system_sysid_qsys_0_control_slave_translator
		generic map (
			AV_ADDRESS_W                   => 1,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 20,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                                               --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                        --                    reset.reset
			uav_address              => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_readdata              => sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_write                 => open,                                                                                  --              (terminated)
			av_read                  => open,                                                                                  --              (terminated)
			av_writedata             => open,                                                                                  --              (terminated)
			av_begintransfer         => open,                                                                                  --              (terminated)
			av_beginbursttransfer    => open,                                                                                  --              (terminated)
			av_burstcount            => open,                                                                                  --              (terminated)
			av_byteenable            => open,                                                                                  --              (terminated)
			av_readdatavalid         => '0',                                                                                   --              (terminated)
			av_waitrequest           => '0',                                                                                   --              (terminated)
			av_writebyteenable       => open,                                                                                  --              (terminated)
			av_lock                  => open,                                                                                  --              (terminated)
			av_chipselect            => open,                                                                                  --              (terminated)
			av_clken                 => open,                                                                                  --              (terminated)
			uav_clken                => '0',                                                                                   --              (terminated)
			av_debugaccess           => open,                                                                                  --              (terminated)
			av_outputenable          => open,                                                                                  --              (terminated)
			uav_response             => open,                                                                                  --              (terminated)
			av_response              => "00",                                                                                  --              (terminated)
			uav_writeresponserequest => '0',                                                                                   --              (terminated)
			uav_writeresponsevalid   => open,                                                                                  --              (terminated)
			av_writeresponserequest  => open,                                                                                  --              (terminated)
			av_writeresponsevalid    => '0'                                                                                    --              (terminated)
		);

	timer_0_s1_translator : component nios_system_timer_0_s1_translator
		generic map (
			AV_ADDRESS_W                   => 3,
			AV_DATA_W                      => 16,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 20,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                               --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                        --                    reset.reset
			uav_address              => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => timer_0_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => timer_0_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => timer_0_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => timer_0_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => timer_0_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                  --              (terminated)
			av_begintransfer         => open,                                                                  --              (terminated)
			av_beginbursttransfer    => open,                                                                  --              (terminated)
			av_burstcount            => open,                                                                  --              (terminated)
			av_byteenable            => open,                                                                  --              (terminated)
			av_readdatavalid         => '0',                                                                   --              (terminated)
			av_waitrequest           => '0',                                                                   --              (terminated)
			av_writebyteenable       => open,                                                                  --              (terminated)
			av_lock                  => open,                                                                  --              (terminated)
			av_clken                 => open,                                                                  --              (terminated)
			uav_clken                => '0',                                                                   --              (terminated)
			av_debugaccess           => open,                                                                  --              (terminated)
			av_outputenable          => open,                                                                  --              (terminated)
			uav_response             => open,                                                                  --              (terminated)
			av_response              => "00",                                                                  --              (terminated)
			uav_writeresponserequest => '0',                                                                   --              (terminated)
			uav_writeresponsevalid   => open,                                                                  --              (terminated)
			av_writeresponserequest  => open,                                                                  --              (terminated)
			av_writeresponsevalid    => '0'                                                                    --              (terminated)
		);

	pio_0_s1_translator : component nios_system_pio_0_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 20,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                             --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                      --                    reset.reset
			uav_address              => pio_0_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => pio_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => pio_0_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => pio_0_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => pio_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => pio_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => pio_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => pio_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => pio_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => pio_0_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => pio_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => pio_0_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => pio_0_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => pio_0_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => pio_0_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => pio_0_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                --              (terminated)
			av_begintransfer         => open,                                                                --              (terminated)
			av_beginbursttransfer    => open,                                                                --              (terminated)
			av_burstcount            => open,                                                                --              (terminated)
			av_byteenable            => open,                                                                --              (terminated)
			av_readdatavalid         => '0',                                                                 --              (terminated)
			av_waitrequest           => '0',                                                                 --              (terminated)
			av_writebyteenable       => open,                                                                --              (terminated)
			av_lock                  => open,                                                                --              (terminated)
			av_clken                 => open,                                                                --              (terminated)
			uav_clken                => '0',                                                                 --              (terminated)
			av_debugaccess           => open,                                                                --              (terminated)
			av_outputenable          => open,                                                                --              (terminated)
			uav_response             => open,                                                                --              (terminated)
			av_response              => "00",                                                                --              (terminated)
			uav_writeresponserequest => '0',                                                                 --              (terminated)
			uav_writeresponsevalid   => open,                                                                --              (terminated)
			av_writeresponserequest  => open,                                                                --              (terminated)
			av_writeresponsevalid    => '0'                                                                  --              (terminated)
		);

	av_status_reg_0_avalon_slave_0_translator : component nios_system_av_status_reg_0_avalon_slave_0_translator
		generic map (
			AV_ADDRESS_W                   => 4,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 20,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                                                   --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                            --                    reset.reset
			uav_address              => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => av_status_reg_0_avalon_slave_0_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => av_status_reg_0_avalon_slave_0_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => av_status_reg_0_avalon_slave_0_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => av_status_reg_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => av_status_reg_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_begintransfer         => open,                                                                                      --              (terminated)
			av_beginbursttransfer    => open,                                                                                      --              (terminated)
			av_burstcount            => open,                                                                                      --              (terminated)
			av_byteenable            => open,                                                                                      --              (terminated)
			av_readdatavalid         => '0',                                                                                       --              (terminated)
			av_waitrequest           => '0',                                                                                       --              (terminated)
			av_writebyteenable       => open,                                                                                      --              (terminated)
			av_lock                  => open,                                                                                      --              (terminated)
			av_chipselect            => open,                                                                                      --              (terminated)
			av_clken                 => open,                                                                                      --              (terminated)
			uav_clken                => '0',                                                                                       --              (terminated)
			av_debugaccess           => open,                                                                                      --              (terminated)
			av_outputenable          => open,                                                                                      --              (terminated)
			uav_response             => open,                                                                                      --              (terminated)
			av_response              => "00",                                                                                      --              (terminated)
			uav_writeresponserequest => '0',                                                                                       --              (terminated)
			uav_writeresponsevalid   => open,                                                                                      --              (terminated)
			av_writeresponserequest  => open,                                                                                      --              (terminated)
			av_writeresponsevalid    => '0'                                                                                        --              (terminated)
		);

	av_eth_config_0_avalon_slave_0_translator : component nios_system_av_status_reg_0_avalon_slave_0_translator
		generic map (
			AV_ADDRESS_W                   => 4,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 20,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                                                   --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                            --                    reset.reset
			uav_address              => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => av_eth_config_0_avalon_slave_0_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => av_eth_config_0_avalon_slave_0_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => av_eth_config_0_avalon_slave_0_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => av_eth_config_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => av_eth_config_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_begintransfer         => open,                                                                                      --              (terminated)
			av_beginbursttransfer    => open,                                                                                      --              (terminated)
			av_burstcount            => open,                                                                                      --              (terminated)
			av_byteenable            => open,                                                                                      --              (terminated)
			av_readdatavalid         => '0',                                                                                       --              (terminated)
			av_waitrequest           => '0',                                                                                       --              (terminated)
			av_writebyteenable       => open,                                                                                      --              (terminated)
			av_lock                  => open,                                                                                      --              (terminated)
			av_chipselect            => open,                                                                                      --              (terminated)
			av_clken                 => open,                                                                                      --              (terminated)
			uav_clken                => '0',                                                                                       --              (terminated)
			av_debugaccess           => open,                                                                                      --              (terminated)
			av_outputenable          => open,                                                                                      --              (terminated)
			uav_response             => open,                                                                                      --              (terminated)
			av_response              => "00",                                                                                      --              (terminated)
			uav_writeresponserequest => '0',                                                                                       --              (terminated)
			uav_writeresponsevalid   => open,                                                                                      --              (terminated)
			av_writeresponserequest  => open,                                                                                      --              (terminated)
			av_writeresponsevalid    => '0'                                                                                        --              (terminated)
		);

	av_config_reg_0_avalon_slave_0_translator : component nios_system_av_status_reg_0_avalon_slave_0_translator
		generic map (
			AV_ADDRESS_W                   => 4,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 20,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                                                   --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                            --                    reset.reset
			uav_address              => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => av_config_reg_0_avalon_slave_0_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => av_config_reg_0_avalon_slave_0_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => av_config_reg_0_avalon_slave_0_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => av_config_reg_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => av_config_reg_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_begintransfer         => open,                                                                                      --              (terminated)
			av_beginbursttransfer    => open,                                                                                      --              (terminated)
			av_burstcount            => open,                                                                                      --              (terminated)
			av_byteenable            => open,                                                                                      --              (terminated)
			av_readdatavalid         => '0',                                                                                       --              (terminated)
			av_waitrequest           => '0',                                                                                       --              (terminated)
			av_writebyteenable       => open,                                                                                      --              (terminated)
			av_lock                  => open,                                                                                      --              (terminated)
			av_chipselect            => open,                                                                                      --              (terminated)
			av_clken                 => open,                                                                                      --              (terminated)
			uav_clken                => '0',                                                                                       --              (terminated)
			av_debugaccess           => open,                                                                                      --              (terminated)
			av_outputenable          => open,                                                                                      --              (terminated)
			uav_response             => open,                                                                                      --              (terminated)
			av_response              => "00",                                                                                      --              (terminated)
			uav_writeresponserequest => '0',                                                                                       --              (terminated)
			uav_writeresponsevalid   => open,                                                                                      --              (terminated)
			av_writeresponserequest  => open,                                                                                      --              (terminated)
			av_writeresponsevalid    => '0'                                                                                        --              (terminated)
		);

	av_sendpacket_0_avalon_slave_0_translator : component nios_system_av_status_reg_0_avalon_slave_0_translator
		generic map (
			AV_ADDRESS_W                   => 4,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 20,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                                                   --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                            --                    reset.reset
			uav_address              => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => av_sendpacket_0_avalon_slave_0_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => av_sendpacket_0_avalon_slave_0_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => av_sendpacket_0_avalon_slave_0_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => av_sendpacket_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => av_sendpacket_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_begintransfer         => open,                                                                                      --              (terminated)
			av_beginbursttransfer    => open,                                                                                      --              (terminated)
			av_burstcount            => open,                                                                                      --              (terminated)
			av_byteenable            => open,                                                                                      --              (terminated)
			av_readdatavalid         => '0',                                                                                       --              (terminated)
			av_waitrequest           => '0',                                                                                       --              (terminated)
			av_writebyteenable       => open,                                                                                      --              (terminated)
			av_lock                  => open,                                                                                      --              (terminated)
			av_chipselect            => open,                                                                                      --              (terminated)
			av_clken                 => open,                                                                                      --              (terminated)
			uav_clken                => '0',                                                                                       --              (terminated)
			av_debugaccess           => open,                                                                                      --              (terminated)
			av_outputenable          => open,                                                                                      --              (terminated)
			uav_response             => open,                                                                                      --              (terminated)
			av_response              => "00",                                                                                      --              (terminated)
			uav_writeresponserequest => '0',                                                                                       --              (terminated)
			uav_writeresponsevalid   => open,                                                                                      --              (terminated)
			av_writeresponserequest  => open,                                                                                      --              (terminated)
			av_writeresponsevalid    => '0'                                                                                        --              (terminated)
		);

	nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent : component altera_merlin_master_agent
		generic map (
			PKT_PROTECTION_H          => 88,
			PKT_PROTECTION_L          => 86,
			PKT_BEGIN_BURST           => 75,
			PKT_BURSTWRAP_H           => 67,
			PKT_BURSTWRAP_L           => 65,
			PKT_BURST_SIZE_H          => 70,
			PKT_BURST_SIZE_L          => 68,
			PKT_BURST_TYPE_H          => 72,
			PKT_BURST_TYPE_L          => 71,
			PKT_BYTE_CNT_H            => 64,
			PKT_BYTE_CNT_L            => 62,
			PKT_ADDR_H                => 55,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 56,
			PKT_TRANS_POSTED          => 57,
			PKT_TRANS_WRITE           => 58,
			PKT_TRANS_READ            => 59,
			PKT_TRANS_LOCK            => 60,
			PKT_TRANS_EXCLUSIVE       => 61,
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_SRC_ID_H              => 80,
			PKT_SRC_ID_L              => 77,
			PKT_DEST_ID_H             => 84,
			PKT_DEST_ID_L             => 81,
			PKT_THREAD_ID_H           => 85,
			PKT_THREAD_ID_L           => 85,
			PKT_CACHE_H               => 92,
			PKT_CACHE_L               => 89,
			PKT_DATA_SIDEBAND_H       => 74,
			PKT_DATA_SIDEBAND_L       => 74,
			PKT_QOS_H                 => 76,
			PKT_QOS_L                 => 76,
			PKT_ADDR_SIDEBAND_H       => 73,
			PKT_ADDR_SIDEBAND_L       => 73,
			PKT_RESPONSE_STATUS_H     => 94,
			PKT_RESPONSE_STATUS_L     => 93,
			ST_DATA_W                 => 95,
			ST_CHANNEL_W              => 10,
			AV_BURSTCOUNT_W           => 3,
			SUPPRESS_0_BYTEEN_RSP     => 0,
			ID                        => 1,
			BURSTWRAP_VALUE           => 3,
			CACHE_VALUE               => 0,
			SECURE_ACCESS_BIT         => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                                     --       clk.clk
			reset                   => rst_controller_reset_out_reset,                                                              -- clk_reset.reset
			av_address              => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_address,                --        av.address
			av_write                => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_write,                  --          .write
			av_read                 => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata            => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata             => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest          => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid        => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable           => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount           => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess          => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock                 => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid                => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data                 => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket        => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket          => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready                => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid                => rsp_xbar_mux_src_valid,                                                                      --        rp.valid
			rp_data                 => rsp_xbar_mux_src_data,                                                                       --          .data
			rp_channel              => rsp_xbar_mux_src_channel,                                                                    --          .channel
			rp_startofpacket        => rsp_xbar_mux_src_startofpacket,                                                              --          .startofpacket
			rp_endofpacket          => rsp_xbar_mux_src_endofpacket,                                                                --          .endofpacket
			rp_ready                => rsp_xbar_mux_src_ready,                                                                      --          .ready
			av_response             => open,                                                                                        -- (terminated)
			av_writeresponserequest => '0',                                                                                         -- (terminated)
			av_writeresponsevalid   => open                                                                                         -- (terminated)
		);

	nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent : component altera_merlin_master_agent
		generic map (
			PKT_PROTECTION_H          => 88,
			PKT_PROTECTION_L          => 86,
			PKT_BEGIN_BURST           => 75,
			PKT_BURSTWRAP_H           => 67,
			PKT_BURSTWRAP_L           => 65,
			PKT_BURST_SIZE_H          => 70,
			PKT_BURST_SIZE_L          => 68,
			PKT_BURST_TYPE_H          => 72,
			PKT_BURST_TYPE_L          => 71,
			PKT_BYTE_CNT_H            => 64,
			PKT_BYTE_CNT_L            => 62,
			PKT_ADDR_H                => 55,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 56,
			PKT_TRANS_POSTED          => 57,
			PKT_TRANS_WRITE           => 58,
			PKT_TRANS_READ            => 59,
			PKT_TRANS_LOCK            => 60,
			PKT_TRANS_EXCLUSIVE       => 61,
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_SRC_ID_H              => 80,
			PKT_SRC_ID_L              => 77,
			PKT_DEST_ID_H             => 84,
			PKT_DEST_ID_L             => 81,
			PKT_THREAD_ID_H           => 85,
			PKT_THREAD_ID_L           => 85,
			PKT_CACHE_H               => 92,
			PKT_CACHE_L               => 89,
			PKT_DATA_SIDEBAND_H       => 74,
			PKT_DATA_SIDEBAND_L       => 74,
			PKT_QOS_H                 => 76,
			PKT_QOS_L                 => 76,
			PKT_ADDR_SIDEBAND_H       => 73,
			PKT_ADDR_SIDEBAND_L       => 73,
			PKT_RESPONSE_STATUS_H     => 94,
			PKT_RESPONSE_STATUS_L     => 93,
			ST_DATA_W                 => 95,
			ST_CHANNEL_W              => 10,
			AV_BURSTCOUNT_W           => 3,
			SUPPRESS_0_BYTEEN_RSP     => 0,
			ID                        => 0,
			BURSTWRAP_VALUE           => 7,
			CACHE_VALUE               => 0,
			SECURE_ACCESS_BIT         => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                              --       clk.clk
			reset                   => rst_controller_reset_out_reset,                                                       -- clk_reset.reset
			av_address              => nios2_qsys_0_data_master_translator_avalon_universal_master_0_address,                --        av.address
			av_write                => nios2_qsys_0_data_master_translator_avalon_universal_master_0_write,                  --          .write
			av_read                 => nios2_qsys_0_data_master_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata            => nios2_qsys_0_data_master_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata             => nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest          => nios2_qsys_0_data_master_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid        => nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable           => nios2_qsys_0_data_master_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount           => nios2_qsys_0_data_master_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess          => nios2_qsys_0_data_master_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock                 => nios2_qsys_0_data_master_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid                => nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data                 => nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket        => nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket          => nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready                => nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid                => rsp_xbar_mux_001_src_valid,                                                           --        rp.valid
			rp_data                 => rsp_xbar_mux_001_src_data,                                                            --          .data
			rp_channel              => rsp_xbar_mux_001_src_channel,                                                         --          .channel
			rp_startofpacket        => rsp_xbar_mux_001_src_startofpacket,                                                   --          .startofpacket
			rp_endofpacket          => rsp_xbar_mux_001_src_endofpacket,                                                     --          .endofpacket
			rp_ready                => rsp_xbar_mux_001_src_ready,                                                           --          .ready
			av_response             => open,                                                                                 -- (terminated)
			av_writeresponserequest => '0',                                                                                  -- (terminated)
			av_writeresponsevalid   => open                                                                                  -- (terminated)
		);

	nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent : component altera_merlin_slave_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 75,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 55,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 56,
			PKT_TRANS_POSTED          => 57,
			PKT_TRANS_WRITE           => 58,
			PKT_TRANS_READ            => 59,
			PKT_TRANS_LOCK            => 60,
			PKT_SRC_ID_H              => 80,
			PKT_SRC_ID_L              => 77,
			PKT_DEST_ID_H             => 84,
			PKT_DEST_ID_L             => 81,
			PKT_BURSTWRAP_H           => 67,
			PKT_BURSTWRAP_L           => 65,
			PKT_BYTE_CNT_H            => 64,
			PKT_BYTE_CNT_L            => 62,
			PKT_PROTECTION_H          => 88,
			PKT_PROTECTION_L          => 86,
			PKT_RESPONSE_STATUS_H     => 94,
			PKT_RESPONSE_STATUS_L     => 93,
			PKT_BURST_SIZE_H          => 70,
			PKT_BURST_SIZE_L          => 68,
			ST_CHANNEL_W              => 10,
			ST_DATA_W                 => 95,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                                             --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                                      --       clk_reset.reset
			m0_address              => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_src_ready,                                                                              --              cp.ready
			cp_valid                => cmd_xbar_mux_src_valid,                                                                              --                .valid
			cp_data                 => cmd_xbar_mux_src_data,                                                                               --                .data
			cp_startofpacket        => cmd_xbar_mux_src_startofpacket,                                                                      --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_src_endofpacket,                                                                        --                .endofpacket
			cp_channel              => cmd_xbar_mux_src_channel,                                                                            --                .channel
			rf_sink_ready           => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                                --     (terminated)
			m0_writeresponserequest => open,                                                                                                --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                                  --     (terminated)
		);

	nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo : component altera_avalon_sc_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 96,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                                             --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                                      -- clk_reset.reset
			in_data           => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                                -- (terminated)
			csr_read          => '0',                                                                                                 -- (terminated)
			csr_write         => '0',                                                                                                 -- (terminated)
			csr_readdata      => open,                                                                                                -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                                  -- (terminated)
			almost_full_data  => open,                                                                                                -- (terminated)
			almost_empty_data => open,                                                                                                -- (terminated)
			in_empty          => '0',                                                                                                 -- (terminated)
			out_empty         => open,                                                                                                -- (terminated)
			in_error          => '0',                                                                                                 -- (terminated)
			out_error         => open,                                                                                                -- (terminated)
			in_channel        => '0',                                                                                                 -- (terminated)
			out_channel       => open                                                                                                 -- (terminated)
		);

	onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent : component altera_merlin_slave_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 75,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 55,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 56,
			PKT_TRANS_POSTED          => 57,
			PKT_TRANS_WRITE           => 58,
			PKT_TRANS_READ            => 59,
			PKT_TRANS_LOCK            => 60,
			PKT_SRC_ID_H              => 80,
			PKT_SRC_ID_L              => 77,
			PKT_DEST_ID_H             => 84,
			PKT_DEST_ID_L             => 81,
			PKT_BURSTWRAP_H           => 67,
			PKT_BURSTWRAP_L           => 65,
			PKT_BYTE_CNT_H            => 64,
			PKT_BYTE_CNT_L            => 62,
			PKT_PROTECTION_H          => 88,
			PKT_PROTECTION_L          => 86,
			PKT_RESPONSE_STATUS_H     => 94,
			PKT_RESPONSE_STATUS_L     => 93,
			PKT_BURST_SIZE_H          => 70,
			PKT_BURST_SIZE_L          => 68,
			ST_CHANNEL_W              => 10,
			ST_DATA_W                 => 95,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                                  --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                           --       clk_reset.reset
			m0_address              => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_001_src_ready,                                                               --              cp.ready
			cp_valid                => cmd_xbar_mux_001_src_valid,                                                               --                .valid
			cp_data                 => cmd_xbar_mux_001_src_data,                                                                --                .data
			cp_startofpacket        => cmd_xbar_mux_001_src_startofpacket,                                                       --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_001_src_endofpacket,                                                         --                .endofpacket
			cp_channel              => cmd_xbar_mux_001_src_channel,                                                             --                .channel
			rf_sink_ready           => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                     --     (terminated)
			m0_writeresponserequest => open,                                                                                     --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                       --     (terminated)
		);

	onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component altera_avalon_sc_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 96,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                                  --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                           -- clk_reset.reset
			in_data           => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                     -- (terminated)
			csr_read          => '0',                                                                                      -- (terminated)
			csr_write         => '0',                                                                                      -- (terminated)
			csr_readdata      => open,                                                                                     -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                       -- (terminated)
			almost_full_data  => open,                                                                                     -- (terminated)
			almost_empty_data => open,                                                                                     -- (terminated)
			in_empty          => '0',                                                                                      -- (terminated)
			out_empty         => open,                                                                                     -- (terminated)
			in_error          => '0',                                                                                      -- (terminated)
			out_error         => open,                                                                                     -- (terminated)
			in_channel        => '0',                                                                                      -- (terminated)
			out_channel       => open                                                                                      -- (terminated)
		);

	jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent : component altera_merlin_slave_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 75,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 55,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 56,
			PKT_TRANS_POSTED          => 57,
			PKT_TRANS_WRITE           => 58,
			PKT_TRANS_READ            => 59,
			PKT_TRANS_LOCK            => 60,
			PKT_SRC_ID_H              => 80,
			PKT_SRC_ID_L              => 77,
			PKT_DEST_ID_H             => 84,
			PKT_DEST_ID_L             => 81,
			PKT_BURSTWRAP_H           => 67,
			PKT_BURSTWRAP_L           => 65,
			PKT_BYTE_CNT_H            => 64,
			PKT_BYTE_CNT_L            => 62,
			PKT_PROTECTION_H          => 88,
			PKT_PROTECTION_L          => 86,
			PKT_RESPONSE_STATUS_H     => 94,
			PKT_RESPONSE_STATUS_L     => 93,
			PKT_BURST_SIZE_H          => 70,
			PKT_BURST_SIZE_L          => 68,
			ST_CHANNEL_W              => 10,
			ST_DATA_W                 => 95,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                                            --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                                     --       clk_reset.reset
			m0_address              => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src2_ready,                                                                      --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src2_valid,                                                                      --                .valid
			cp_data                 => cmd_xbar_demux_001_src2_data,                                                                       --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src2_startofpacket,                                                              --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src2_endofpacket,                                                                --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src2_channel,                                                                    --                .channel
			rf_sink_ready           => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                               --     (terminated)
			m0_writeresponserequest => open,                                                                                               --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                                 --     (terminated)
		);

	jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component altera_avalon_sc_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 96,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                                            --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                                     -- clk_reset.reset
			in_data           => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                               -- (terminated)
			csr_read          => '0',                                                                                                -- (terminated)
			csr_write         => '0',                                                                                                -- (terminated)
			csr_readdata      => open,                                                                                               -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                                 -- (terminated)
			almost_full_data  => open,                                                                                               -- (terminated)
			almost_empty_data => open,                                                                                               -- (terminated)
			in_empty          => '0',                                                                                                -- (terminated)
			out_empty         => open,                                                                                               -- (terminated)
			in_error          => '0',                                                                                                -- (terminated)
			out_error         => open,                                                                                               -- (terminated)
			in_channel        => '0',                                                                                                -- (terminated)
			out_channel       => open                                                                                                -- (terminated)
		);

	sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent : component altera_merlin_slave_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 75,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 55,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 56,
			PKT_TRANS_POSTED          => 57,
			PKT_TRANS_WRITE           => 58,
			PKT_TRANS_READ            => 59,
			PKT_TRANS_LOCK            => 60,
			PKT_SRC_ID_H              => 80,
			PKT_SRC_ID_L              => 77,
			PKT_DEST_ID_H             => 84,
			PKT_DEST_ID_L             => 81,
			PKT_BURSTWRAP_H           => 67,
			PKT_BURSTWRAP_L           => 65,
			PKT_BYTE_CNT_H            => 64,
			PKT_BYTE_CNT_L            => 62,
			PKT_PROTECTION_H          => 88,
			PKT_PROTECTION_L          => 86,
			PKT_RESPONSE_STATUS_H     => 94,
			PKT_RESPONSE_STATUS_L     => 93,
			PKT_BURST_SIZE_H          => 70,
			PKT_BURST_SIZE_L          => 68,
			ST_CHANNEL_W              => 10,
			ST_DATA_W                 => 95,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                                         --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                                  --       clk_reset.reset
			m0_address              => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src3_ready,                                                                   --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src3_valid,                                                                   --                .valid
			cp_data                 => cmd_xbar_demux_001_src3_data,                                                                    --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src3_startofpacket,                                                           --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src3_endofpacket,                                                             --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src3_channel,                                                                 --                .channel
			rf_sink_ready           => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                            --     (terminated)
			m0_writeresponserequest => open,                                                                                            --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                              --     (terminated)
		);

	sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component altera_avalon_sc_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 96,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                                         --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                                  -- clk_reset.reset
			in_data           => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                            -- (terminated)
			csr_read          => '0',                                                                                             -- (terminated)
			csr_write         => '0',                                                                                             -- (terminated)
			csr_readdata      => open,                                                                                            -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                              -- (terminated)
			almost_full_data  => open,                                                                                            -- (terminated)
			almost_empty_data => open,                                                                                            -- (terminated)
			in_empty          => '0',                                                                                             -- (terminated)
			out_empty         => open,                                                                                            -- (terminated)
			in_error          => '0',                                                                                             -- (terminated)
			out_error         => open,                                                                                            -- (terminated)
			in_channel        => '0',                                                                                             -- (terminated)
			out_channel       => open                                                                                             -- (terminated)
		);

	timer_0_s1_translator_avalon_universal_slave_0_agent : component altera_merlin_slave_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 75,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 55,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 56,
			PKT_TRANS_POSTED          => 57,
			PKT_TRANS_WRITE           => 58,
			PKT_TRANS_READ            => 59,
			PKT_TRANS_LOCK            => 60,
			PKT_SRC_ID_H              => 80,
			PKT_SRC_ID_L              => 77,
			PKT_DEST_ID_H             => 84,
			PKT_DEST_ID_L             => 81,
			PKT_BURSTWRAP_H           => 67,
			PKT_BURSTWRAP_L           => 65,
			PKT_BYTE_CNT_H            => 64,
			PKT_BYTE_CNT_L            => 62,
			PKT_PROTECTION_H          => 88,
			PKT_PROTECTION_L          => 86,
			PKT_RESPONSE_STATUS_H     => 94,
			PKT_RESPONSE_STATUS_L     => 93,
			PKT_BURST_SIZE_H          => 70,
			PKT_BURST_SIZE_L          => 68,
			ST_CHANNEL_W              => 10,
			ST_DATA_W                 => 95,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                         --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                  --       clk_reset.reset
			m0_address              => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src4_ready,                                                   --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src4_valid,                                                   --                .valid
			cp_data                 => cmd_xbar_demux_001_src4_data,                                                    --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src4_startofpacket,                                           --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src4_endofpacket,                                             --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src4_channel,                                                 --                .channel
			rf_sink_ready           => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                            --     (terminated)
			m0_writeresponserequest => open,                                                                            --     (terminated)
			m0_writeresponsevalid   => '0'                                                                              --     (terminated)
		);

	timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component altera_avalon_sc_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 96,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                         --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                  -- clk_reset.reset
			in_data           => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                            -- (terminated)
			csr_read          => '0',                                                                             -- (terminated)
			csr_write         => '0',                                                                             -- (terminated)
			csr_readdata      => open,                                                                            -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                              -- (terminated)
			almost_full_data  => open,                                                                            -- (terminated)
			almost_empty_data => open,                                                                            -- (terminated)
			in_empty          => '0',                                                                             -- (terminated)
			out_empty         => open,                                                                            -- (terminated)
			in_error          => '0',                                                                             -- (terminated)
			out_error         => open,                                                                            -- (terminated)
			in_channel        => '0',                                                                             -- (terminated)
			out_channel       => open                                                                             -- (terminated)
		);

	pio_0_s1_translator_avalon_universal_slave_0_agent : component altera_merlin_slave_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 75,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 55,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 56,
			PKT_TRANS_POSTED          => 57,
			PKT_TRANS_WRITE           => 58,
			PKT_TRANS_READ            => 59,
			PKT_TRANS_LOCK            => 60,
			PKT_SRC_ID_H              => 80,
			PKT_SRC_ID_L              => 77,
			PKT_DEST_ID_H             => 84,
			PKT_DEST_ID_L             => 81,
			PKT_BURSTWRAP_H           => 67,
			PKT_BURSTWRAP_L           => 65,
			PKT_BYTE_CNT_H            => 64,
			PKT_BYTE_CNT_L            => 62,
			PKT_PROTECTION_H          => 88,
			PKT_PROTECTION_L          => 86,
			PKT_RESPONSE_STATUS_H     => 94,
			PKT_RESPONSE_STATUS_L     => 93,
			PKT_BURST_SIZE_H          => 70,
			PKT_BURST_SIZE_L          => 68,
			ST_CHANNEL_W              => 10,
			ST_DATA_W                 => 95,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                       --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                --       clk_reset.reset
			m0_address              => pio_0_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => pio_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => pio_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => pio_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => pio_0_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => pio_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => pio_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => pio_0_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => pio_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => pio_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => pio_0_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => pio_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => pio_0_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => pio_0_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => pio_0_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => pio_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src5_ready,                                                 --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src5_valid,                                                 --                .valid
			cp_data                 => cmd_xbar_demux_001_src5_data,                                                  --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src5_startofpacket,                                         --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src5_endofpacket,                                           --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src5_channel,                                               --                .channel
			rf_sink_ready           => pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                          --     (terminated)
			m0_writeresponserequest => open,                                                                          --     (terminated)
			m0_writeresponsevalid   => '0'                                                                            --     (terminated)
		);

	pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component altera_avalon_sc_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 96,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                       --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                -- clk_reset.reset
			in_data           => pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                          -- (terminated)
			csr_read          => '0',                                                                           -- (terminated)
			csr_write         => '0',                                                                           -- (terminated)
			csr_readdata      => open,                                                                          -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                            -- (terminated)
			almost_full_data  => open,                                                                          -- (terminated)
			almost_empty_data => open,                                                                          -- (terminated)
			in_empty          => '0',                                                                           -- (terminated)
			out_empty         => open,                                                                          -- (terminated)
			in_error          => '0',                                                                           -- (terminated)
			out_error         => open,                                                                          -- (terminated)
			in_channel        => '0',                                                                           -- (terminated)
			out_channel       => open                                                                           -- (terminated)
		);

	av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent : component altera_merlin_slave_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 75,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 55,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 56,
			PKT_TRANS_POSTED          => 57,
			PKT_TRANS_WRITE           => 58,
			PKT_TRANS_READ            => 59,
			PKT_TRANS_LOCK            => 60,
			PKT_SRC_ID_H              => 80,
			PKT_SRC_ID_L              => 77,
			PKT_DEST_ID_H             => 84,
			PKT_DEST_ID_L             => 81,
			PKT_BURSTWRAP_H           => 67,
			PKT_BURSTWRAP_L           => 65,
			PKT_BYTE_CNT_H            => 64,
			PKT_BYTE_CNT_L            => 62,
			PKT_PROTECTION_H          => 88,
			PKT_PROTECTION_L          => 86,
			PKT_RESPONSE_STATUS_H     => 94,
			PKT_RESPONSE_STATUS_L     => 93,
			PKT_BURST_SIZE_H          => 70,
			PKT_BURST_SIZE_L          => 68,
			ST_CHANNEL_W              => 10,
			ST_DATA_W                 => 95,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                                             --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                                      --       clk_reset.reset
			m0_address              => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src6_ready,                                                                       --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src6_valid,                                                                       --                .valid
			cp_data                 => cmd_xbar_demux_001_src6_data,                                                                        --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src6_startofpacket,                                                               --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src6_endofpacket,                                                                 --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src6_channel,                                                                     --                .channel
			rf_sink_ready           => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                                --     (terminated)
			m0_writeresponserequest => open,                                                                                                --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                                  --     (terminated)
		);

	av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo : component altera_avalon_sc_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 96,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                                             --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                                      -- clk_reset.reset
			in_data           => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                                -- (terminated)
			csr_read          => '0',                                                                                                 -- (terminated)
			csr_write         => '0',                                                                                                 -- (terminated)
			csr_readdata      => open,                                                                                                -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                                  -- (terminated)
			almost_full_data  => open,                                                                                                -- (terminated)
			almost_empty_data => open,                                                                                                -- (terminated)
			in_empty          => '0',                                                                                                 -- (terminated)
			out_empty         => open,                                                                                                -- (terminated)
			in_error          => '0',                                                                                                 -- (terminated)
			out_error         => open,                                                                                                -- (terminated)
			in_channel        => '0',                                                                                                 -- (terminated)
			out_channel       => open                                                                                                 -- (terminated)
		);

	av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent : component altera_merlin_slave_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 75,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 55,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 56,
			PKT_TRANS_POSTED          => 57,
			PKT_TRANS_WRITE           => 58,
			PKT_TRANS_READ            => 59,
			PKT_TRANS_LOCK            => 60,
			PKT_SRC_ID_H              => 80,
			PKT_SRC_ID_L              => 77,
			PKT_DEST_ID_H             => 84,
			PKT_DEST_ID_L             => 81,
			PKT_BURSTWRAP_H           => 67,
			PKT_BURSTWRAP_L           => 65,
			PKT_BYTE_CNT_H            => 64,
			PKT_BYTE_CNT_L            => 62,
			PKT_PROTECTION_H          => 88,
			PKT_PROTECTION_L          => 86,
			PKT_RESPONSE_STATUS_H     => 94,
			PKT_RESPONSE_STATUS_L     => 93,
			PKT_BURST_SIZE_H          => 70,
			PKT_BURST_SIZE_L          => 68,
			ST_CHANNEL_W              => 10,
			ST_DATA_W                 => 95,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                                             --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                                      --       clk_reset.reset
			m0_address              => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src7_ready,                                                                       --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src7_valid,                                                                       --                .valid
			cp_data                 => cmd_xbar_demux_001_src7_data,                                                                        --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src7_startofpacket,                                                               --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src7_endofpacket,                                                                 --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src7_channel,                                                                     --                .channel
			rf_sink_ready           => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                                --     (terminated)
			m0_writeresponserequest => open,                                                                                                --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                                  --     (terminated)
		);

	av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo : component altera_avalon_sc_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 96,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                                             --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                                      -- clk_reset.reset
			in_data           => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                                -- (terminated)
			csr_read          => '0',                                                                                                 -- (terminated)
			csr_write         => '0',                                                                                                 -- (terminated)
			csr_readdata      => open,                                                                                                -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                                  -- (terminated)
			almost_full_data  => open,                                                                                                -- (terminated)
			almost_empty_data => open,                                                                                                -- (terminated)
			in_empty          => '0',                                                                                                 -- (terminated)
			out_empty         => open,                                                                                                -- (terminated)
			in_error          => '0',                                                                                                 -- (terminated)
			out_error         => open,                                                                                                -- (terminated)
			in_channel        => '0',                                                                                                 -- (terminated)
			out_channel       => open                                                                                                 -- (terminated)
		);

	av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent : component altera_merlin_slave_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 75,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 55,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 56,
			PKT_TRANS_POSTED          => 57,
			PKT_TRANS_WRITE           => 58,
			PKT_TRANS_READ            => 59,
			PKT_TRANS_LOCK            => 60,
			PKT_SRC_ID_H              => 80,
			PKT_SRC_ID_L              => 77,
			PKT_DEST_ID_H             => 84,
			PKT_DEST_ID_L             => 81,
			PKT_BURSTWRAP_H           => 67,
			PKT_BURSTWRAP_L           => 65,
			PKT_BYTE_CNT_H            => 64,
			PKT_BYTE_CNT_L            => 62,
			PKT_PROTECTION_H          => 88,
			PKT_PROTECTION_L          => 86,
			PKT_RESPONSE_STATUS_H     => 94,
			PKT_RESPONSE_STATUS_L     => 93,
			PKT_BURST_SIZE_H          => 70,
			PKT_BURST_SIZE_L          => 68,
			ST_CHANNEL_W              => 10,
			ST_DATA_W                 => 95,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                                             --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                                      --       clk_reset.reset
			m0_address              => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src8_ready,                                                                       --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src8_valid,                                                                       --                .valid
			cp_data                 => cmd_xbar_demux_001_src8_data,                                                                        --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src8_startofpacket,                                                               --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src8_endofpacket,                                                                 --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src8_channel,                                                                     --                .channel
			rf_sink_ready           => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                                --     (terminated)
			m0_writeresponserequest => open,                                                                                                --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                                  --     (terminated)
		);

	av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo : component altera_avalon_sc_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 96,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                                             --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                                      -- clk_reset.reset
			in_data           => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                                -- (terminated)
			csr_read          => '0',                                                                                                 -- (terminated)
			csr_write         => '0',                                                                                                 -- (terminated)
			csr_readdata      => open,                                                                                                -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                                  -- (terminated)
			almost_full_data  => open,                                                                                                -- (terminated)
			almost_empty_data => open,                                                                                                -- (terminated)
			in_empty          => '0',                                                                                                 -- (terminated)
			out_empty         => open,                                                                                                -- (terminated)
			in_error          => '0',                                                                                                 -- (terminated)
			out_error         => open,                                                                                                -- (terminated)
			in_channel        => '0',                                                                                                 -- (terminated)
			out_channel       => open                                                                                                 -- (terminated)
		);

	av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent : component altera_merlin_slave_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 75,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 55,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 56,
			PKT_TRANS_POSTED          => 57,
			PKT_TRANS_WRITE           => 58,
			PKT_TRANS_READ            => 59,
			PKT_TRANS_LOCK            => 60,
			PKT_SRC_ID_H              => 80,
			PKT_SRC_ID_L              => 77,
			PKT_DEST_ID_H             => 84,
			PKT_DEST_ID_L             => 81,
			PKT_BURSTWRAP_H           => 67,
			PKT_BURSTWRAP_L           => 65,
			PKT_BYTE_CNT_H            => 64,
			PKT_BYTE_CNT_L            => 62,
			PKT_PROTECTION_H          => 88,
			PKT_PROTECTION_L          => 86,
			PKT_RESPONSE_STATUS_H     => 94,
			PKT_RESPONSE_STATUS_L     => 93,
			PKT_BURST_SIZE_H          => 70,
			PKT_BURST_SIZE_L          => 68,
			ST_CHANNEL_W              => 10,
			ST_DATA_W                 => 95,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                                             --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                                      --       clk_reset.reset
			m0_address              => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src9_ready,                                                                       --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src9_valid,                                                                       --                .valid
			cp_data                 => cmd_xbar_demux_001_src9_data,                                                                        --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src9_startofpacket,                                                               --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src9_endofpacket,                                                                 --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src9_channel,                                                                     --                .channel
			rf_sink_ready           => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                                --     (terminated)
			m0_writeresponserequest => open,                                                                                                --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                                  --     (terminated)
		);

	av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo : component altera_avalon_sc_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 96,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                                             --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                                      -- clk_reset.reset
			in_data           => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                                -- (terminated)
			csr_read          => '0',                                                                                                 -- (terminated)
			csr_write         => '0',                                                                                                 -- (terminated)
			csr_readdata      => open,                                                                                                -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                                  -- (terminated)
			almost_full_data  => open,                                                                                                -- (terminated)
			almost_empty_data => open,                                                                                                -- (terminated)
			in_empty          => '0',                                                                                                 -- (terminated)
			out_empty         => open,                                                                                                -- (terminated)
			in_error          => '0',                                                                                                 -- (terminated)
			out_error         => open,                                                                                                -- (terminated)
			in_channel        => '0',                                                                                                 -- (terminated)
			out_channel       => open                                                                                                 -- (terminated)
		);

	addr_router : component nios_system_addr_router
		port map (
			sink_ready         => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                                     --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                              -- clk_reset.reset
			src_ready          => addr_router_src_ready,                                                                       --       src.ready
			src_valid          => addr_router_src_valid,                                                                       --          .valid
			src_data           => addr_router_src_data,                                                                        --          .data
			src_channel        => addr_router_src_channel,                                                                     --          .channel
			src_startofpacket  => addr_router_src_startofpacket,                                                               --          .startofpacket
			src_endofpacket    => addr_router_src_endofpacket                                                                  --          .endofpacket
		);

	addr_router_001 : component nios_system_addr_router_001
		port map (
			sink_ready         => nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                              --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                       -- clk_reset.reset
			src_ready          => addr_router_001_src_ready,                                                            --       src.ready
			src_valid          => addr_router_001_src_valid,                                                            --          .valid
			src_data           => addr_router_001_src_data,                                                             --          .data
			src_channel        => addr_router_001_src_channel,                                                          --          .channel
			src_startofpacket  => addr_router_001_src_startofpacket,                                                    --          .startofpacket
			src_endofpacket    => addr_router_001_src_endofpacket                                                       --          .endofpacket
		);

	id_router : component nios_system_id_router
		port map (
			sink_ready         => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                                   --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                            -- clk_reset.reset
			src_ready          => id_router_src_ready,                                                                       --       src.ready
			src_valid          => id_router_src_valid,                                                                       --          .valid
			src_data           => id_router_src_data,                                                                        --          .data
			src_channel        => id_router_src_channel,                                                                     --          .channel
			src_startofpacket  => id_router_src_startofpacket,                                                               --          .startofpacket
			src_endofpacket    => id_router_src_endofpacket                                                                  --          .endofpacket
		);

	id_router_001 : component nios_system_id_router
		port map (
			sink_ready         => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                        --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                 -- clk_reset.reset
			src_ready          => id_router_001_src_ready,                                                        --       src.ready
			src_valid          => id_router_001_src_valid,                                                        --          .valid
			src_data           => id_router_001_src_data,                                                         --          .data
			src_channel        => id_router_001_src_channel,                                                      --          .channel
			src_startofpacket  => id_router_001_src_startofpacket,                                                --          .startofpacket
			src_endofpacket    => id_router_001_src_endofpacket                                                   --          .endofpacket
		);

	id_router_002 : component nios_system_id_router_002
		port map (
			sink_ready         => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                                  --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                           -- clk_reset.reset
			src_ready          => id_router_002_src_ready,                                                                  --       src.ready
			src_valid          => id_router_002_src_valid,                                                                  --          .valid
			src_data           => id_router_002_src_data,                                                                   --          .data
			src_channel        => id_router_002_src_channel,                                                                --          .channel
			src_startofpacket  => id_router_002_src_startofpacket,                                                          --          .startofpacket
			src_endofpacket    => id_router_002_src_endofpacket                                                             --          .endofpacket
		);

	id_router_003 : component nios_system_id_router_002
		port map (
			sink_ready         => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                               --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                        -- clk_reset.reset
			src_ready          => id_router_003_src_ready,                                                               --       src.ready
			src_valid          => id_router_003_src_valid,                                                               --          .valid
			src_data           => id_router_003_src_data,                                                                --          .data
			src_channel        => id_router_003_src_channel,                                                             --          .channel
			src_startofpacket  => id_router_003_src_startofpacket,                                                       --          .startofpacket
			src_endofpacket    => id_router_003_src_endofpacket                                                          --          .endofpacket
		);

	id_router_004 : component nios_system_id_router_002
		port map (
			sink_ready         => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                               --       clk.clk
			reset              => rst_controller_reset_out_reset,                                        -- clk_reset.reset
			src_ready          => id_router_004_src_ready,                                               --       src.ready
			src_valid          => id_router_004_src_valid,                                               --          .valid
			src_data           => id_router_004_src_data,                                                --          .data
			src_channel        => id_router_004_src_channel,                                             --          .channel
			src_startofpacket  => id_router_004_src_startofpacket,                                       --          .startofpacket
			src_endofpacket    => id_router_004_src_endofpacket                                          --          .endofpacket
		);

	id_router_005 : component nios_system_id_router_002
		port map (
			sink_ready         => pio_0_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => pio_0_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => pio_0_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => pio_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => pio_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                             --       clk.clk
			reset              => rst_controller_reset_out_reset,                                      -- clk_reset.reset
			src_ready          => id_router_005_src_ready,                                             --       src.ready
			src_valid          => id_router_005_src_valid,                                             --          .valid
			src_data           => id_router_005_src_data,                                              --          .data
			src_channel        => id_router_005_src_channel,                                           --          .channel
			src_startofpacket  => id_router_005_src_startofpacket,                                     --          .startofpacket
			src_endofpacket    => id_router_005_src_endofpacket                                        --          .endofpacket
		);

	id_router_006 : component nios_system_id_router_002
		port map (
			sink_ready         => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => av_status_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                                   --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                            -- clk_reset.reset
			src_ready          => id_router_006_src_ready,                                                                   --       src.ready
			src_valid          => id_router_006_src_valid,                                                                   --          .valid
			src_data           => id_router_006_src_data,                                                                    --          .data
			src_channel        => id_router_006_src_channel,                                                                 --          .channel
			src_startofpacket  => id_router_006_src_startofpacket,                                                           --          .startofpacket
			src_endofpacket    => id_router_006_src_endofpacket                                                              --          .endofpacket
		);

	id_router_007 : component nios_system_id_router_002
		port map (
			sink_ready         => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => av_eth_config_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                                   --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                            -- clk_reset.reset
			src_ready          => id_router_007_src_ready,                                                                   --       src.ready
			src_valid          => id_router_007_src_valid,                                                                   --          .valid
			src_data           => id_router_007_src_data,                                                                    --          .data
			src_channel        => id_router_007_src_channel,                                                                 --          .channel
			src_startofpacket  => id_router_007_src_startofpacket,                                                           --          .startofpacket
			src_endofpacket    => id_router_007_src_endofpacket                                                              --          .endofpacket
		);

	id_router_008 : component nios_system_id_router_002
		port map (
			sink_ready         => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => av_config_reg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                                   --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                            -- clk_reset.reset
			src_ready          => id_router_008_src_ready,                                                                   --       src.ready
			src_valid          => id_router_008_src_valid,                                                                   --          .valid
			src_data           => id_router_008_src_data,                                                                    --          .data
			src_channel        => id_router_008_src_channel,                                                                 --          .channel
			src_startofpacket  => id_router_008_src_startofpacket,                                                           --          .startofpacket
			src_endofpacket    => id_router_008_src_endofpacket                                                              --          .endofpacket
		);

	id_router_009 : component nios_system_id_router_002
		port map (
			sink_ready         => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => av_sendpacket_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                                   --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                            -- clk_reset.reset
			src_ready          => id_router_009_src_ready,                                                                   --       src.ready
			src_valid          => id_router_009_src_valid,                                                                   --          .valid
			src_data           => id_router_009_src_data,                                                                    --          .data
			src_channel        => id_router_009_src_channel,                                                                 --          .channel
			src_startofpacket  => id_router_009_src_startofpacket,                                                           --          .startofpacket
			src_endofpacket    => id_router_009_src_endofpacket                                                              --          .endofpacket
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS        => 1,
			OUTPUT_RESET_SYNC_EDGES => "deassert",
			SYNC_DEPTH              => 2
		)
		port map (
			reset_in0  => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk        => clk_clk,                        --       clk.clk
			reset_out  => rst_controller_reset_out_reset, -- reset_out.reset
			reset_in1  => '0',                            -- (terminated)
			reset_in2  => '0',                            -- (terminated)
			reset_in3  => '0',                            -- (terminated)
			reset_in4  => '0',                            -- (terminated)
			reset_in5  => '0',                            -- (terminated)
			reset_in6  => '0',                            -- (terminated)
			reset_in7  => '0',                            -- (terminated)
			reset_in8  => '0',                            -- (terminated)
			reset_in9  => '0',                            -- (terminated)
			reset_in10 => '0',                            -- (terminated)
			reset_in11 => '0',                            -- (terminated)
			reset_in12 => '0',                            -- (terminated)
			reset_in13 => '0',                            -- (terminated)
			reset_in14 => '0',                            -- (terminated)
			reset_in15 => '0'                             -- (terminated)
		);

	cmd_xbar_demux : component nios_system_cmd_xbar_demux
		port map (
			clk                => clk_clk,                           --       clk.clk
			reset              => rst_controller_reset_out_reset,    -- clk_reset.reset
			sink_ready         => addr_router_src_ready,             --      sink.ready
			sink_channel       => addr_router_src_channel,           --          .channel
			sink_data          => addr_router_src_data,              --          .data
			sink_startofpacket => addr_router_src_startofpacket,     --          .startofpacket
			sink_endofpacket   => addr_router_src_endofpacket,       --          .endofpacket
			sink_valid(0)      => addr_router_src_valid,             --          .valid
			src0_ready         => cmd_xbar_demux_src0_ready,         --      src0.ready
			src0_valid         => cmd_xbar_demux_src0_valid,         --          .valid
			src0_data          => cmd_xbar_demux_src0_data,          --          .data
			src0_channel       => cmd_xbar_demux_src0_channel,       --          .channel
			src0_startofpacket => cmd_xbar_demux_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => cmd_xbar_demux_src0_endofpacket,   --          .endofpacket
			src1_ready         => cmd_xbar_demux_src1_ready,         --      src1.ready
			src1_valid         => cmd_xbar_demux_src1_valid,         --          .valid
			src1_data          => cmd_xbar_demux_src1_data,          --          .data
			src1_channel       => cmd_xbar_demux_src1_channel,       --          .channel
			src1_startofpacket => cmd_xbar_demux_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => cmd_xbar_demux_src1_endofpacket    --          .endofpacket
		);

	cmd_xbar_demux_001 : component nios_system_cmd_xbar_demux_001
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => addr_router_001_src_ready,             --      sink.ready
			sink_channel       => addr_router_001_src_channel,           --          .channel
			sink_data          => addr_router_001_src_data,              --          .data
			sink_startofpacket => addr_router_001_src_startofpacket,     --          .startofpacket
			sink_endofpacket   => addr_router_001_src_endofpacket,       --          .endofpacket
			sink_valid(0)      => addr_router_001_src_valid,             --          .valid
			src0_ready         => cmd_xbar_demux_001_src0_ready,         --      src0.ready
			src0_valid         => cmd_xbar_demux_001_src0_valid,         --          .valid
			src0_data          => cmd_xbar_demux_001_src0_data,          --          .data
			src0_channel       => cmd_xbar_demux_001_src0_channel,       --          .channel
			src0_startofpacket => cmd_xbar_demux_001_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => cmd_xbar_demux_001_src0_endofpacket,   --          .endofpacket
			src1_ready         => cmd_xbar_demux_001_src1_ready,         --      src1.ready
			src1_valid         => cmd_xbar_demux_001_src1_valid,         --          .valid
			src1_data          => cmd_xbar_demux_001_src1_data,          --          .data
			src1_channel       => cmd_xbar_demux_001_src1_channel,       --          .channel
			src1_startofpacket => cmd_xbar_demux_001_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => cmd_xbar_demux_001_src1_endofpacket,   --          .endofpacket
			src2_ready         => cmd_xbar_demux_001_src2_ready,         --      src2.ready
			src2_valid         => cmd_xbar_demux_001_src2_valid,         --          .valid
			src2_data          => cmd_xbar_demux_001_src2_data,          --          .data
			src2_channel       => cmd_xbar_demux_001_src2_channel,       --          .channel
			src2_startofpacket => cmd_xbar_demux_001_src2_startofpacket, --          .startofpacket
			src2_endofpacket   => cmd_xbar_demux_001_src2_endofpacket,   --          .endofpacket
			src3_ready         => cmd_xbar_demux_001_src3_ready,         --      src3.ready
			src3_valid         => cmd_xbar_demux_001_src3_valid,         --          .valid
			src3_data          => cmd_xbar_demux_001_src3_data,          --          .data
			src3_channel       => cmd_xbar_demux_001_src3_channel,       --          .channel
			src3_startofpacket => cmd_xbar_demux_001_src3_startofpacket, --          .startofpacket
			src3_endofpacket   => cmd_xbar_demux_001_src3_endofpacket,   --          .endofpacket
			src4_ready         => cmd_xbar_demux_001_src4_ready,         --      src4.ready
			src4_valid         => cmd_xbar_demux_001_src4_valid,         --          .valid
			src4_data          => cmd_xbar_demux_001_src4_data,          --          .data
			src4_channel       => cmd_xbar_demux_001_src4_channel,       --          .channel
			src4_startofpacket => cmd_xbar_demux_001_src4_startofpacket, --          .startofpacket
			src4_endofpacket   => cmd_xbar_demux_001_src4_endofpacket,   --          .endofpacket
			src5_ready         => cmd_xbar_demux_001_src5_ready,         --      src5.ready
			src5_valid         => cmd_xbar_demux_001_src5_valid,         --          .valid
			src5_data          => cmd_xbar_demux_001_src5_data,          --          .data
			src5_channel       => cmd_xbar_demux_001_src5_channel,       --          .channel
			src5_startofpacket => cmd_xbar_demux_001_src5_startofpacket, --          .startofpacket
			src5_endofpacket   => cmd_xbar_demux_001_src5_endofpacket,   --          .endofpacket
			src6_ready         => cmd_xbar_demux_001_src6_ready,         --      src6.ready
			src6_valid         => cmd_xbar_demux_001_src6_valid,         --          .valid
			src6_data          => cmd_xbar_demux_001_src6_data,          --          .data
			src6_channel       => cmd_xbar_demux_001_src6_channel,       --          .channel
			src6_startofpacket => cmd_xbar_demux_001_src6_startofpacket, --          .startofpacket
			src6_endofpacket   => cmd_xbar_demux_001_src6_endofpacket,   --          .endofpacket
			src7_ready         => cmd_xbar_demux_001_src7_ready,         --      src7.ready
			src7_valid         => cmd_xbar_demux_001_src7_valid,         --          .valid
			src7_data          => cmd_xbar_demux_001_src7_data,          --          .data
			src7_channel       => cmd_xbar_demux_001_src7_channel,       --          .channel
			src7_startofpacket => cmd_xbar_demux_001_src7_startofpacket, --          .startofpacket
			src7_endofpacket   => cmd_xbar_demux_001_src7_endofpacket,   --          .endofpacket
			src8_ready         => cmd_xbar_demux_001_src8_ready,         --      src8.ready
			src8_valid         => cmd_xbar_demux_001_src8_valid,         --          .valid
			src8_data          => cmd_xbar_demux_001_src8_data,          --          .data
			src8_channel       => cmd_xbar_demux_001_src8_channel,       --          .channel
			src8_startofpacket => cmd_xbar_demux_001_src8_startofpacket, --          .startofpacket
			src8_endofpacket   => cmd_xbar_demux_001_src8_endofpacket,   --          .endofpacket
			src9_ready         => cmd_xbar_demux_001_src9_ready,         --      src9.ready
			src9_valid         => cmd_xbar_demux_001_src9_valid,         --          .valid
			src9_data          => cmd_xbar_demux_001_src9_data,          --          .data
			src9_channel       => cmd_xbar_demux_001_src9_channel,       --          .channel
			src9_startofpacket => cmd_xbar_demux_001_src9_startofpacket, --          .startofpacket
			src9_endofpacket   => cmd_xbar_demux_001_src9_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux : component nios_system_cmd_xbar_mux
		port map (
			clk                 => clk_clk,                               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_src_ready,                --       src.ready
			src_valid           => cmd_xbar_mux_src_valid,                --          .valid
			src_data            => cmd_xbar_mux_src_data,                 --          .data
			src_channel         => cmd_xbar_mux_src_channel,              --          .channel
			src_startofpacket   => cmd_xbar_mux_src_startofpacket,        --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_src_endofpacket,          --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src0_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src0_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src0_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src0_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src0_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src0_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src0_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src0_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src0_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src0_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src0_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src0_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_001 : component nios_system_cmd_xbar_mux
		port map (
			clk                 => clk_clk,                               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_001_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_001_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_001_src_data,             --          .data
			src_channel         => cmd_xbar_mux_001_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_001_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_001_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src1_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src1_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src1_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src1_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src1_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src1_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src1_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src1_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src1_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src1_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src1_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux : component nios_system_cmd_xbar_demux
		port map (
			clk                => clk_clk,                           --       clk.clk
			reset              => rst_controller_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_src_ready,               --      sink.ready
			sink_channel       => id_router_src_channel,             --          .channel
			sink_data          => id_router_src_data,                --          .data
			sink_startofpacket => id_router_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_001 : component nios_system_cmd_xbar_demux
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_001_src_ready,               --      sink.ready
			sink_channel       => id_router_001_src_channel,             --          .channel
			sink_data          => id_router_001_src_data,                --          .data
			sink_startofpacket => id_router_001_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_001_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_001_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_001_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_001_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_001_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_001_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_001_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_001_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_001_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_001_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_001_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_001_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_001_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_001_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_002 : component nios_system_rsp_xbar_demux_002
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_002_src_ready,               --      sink.ready
			sink_channel       => id_router_002_src_channel,             --          .channel
			sink_data          => id_router_002_src_data,                --          .data
			sink_startofpacket => id_router_002_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_002_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_002_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_002_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_002_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_002_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_002_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_002_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_002_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_003 : component nios_system_rsp_xbar_demux_002
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_003_src_ready,               --      sink.ready
			sink_channel       => id_router_003_src_channel,             --          .channel
			sink_data          => id_router_003_src_data,                --          .data
			sink_startofpacket => id_router_003_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_003_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_003_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_003_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_003_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_003_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_003_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_003_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_003_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_004 : component nios_system_rsp_xbar_demux_002
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_004_src_ready,               --      sink.ready
			sink_channel       => id_router_004_src_channel,             --          .channel
			sink_data          => id_router_004_src_data,                --          .data
			sink_startofpacket => id_router_004_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_004_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_004_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_004_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_004_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_004_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_004_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_004_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_004_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_005 : component nios_system_rsp_xbar_demux_002
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_005_src_ready,               --      sink.ready
			sink_channel       => id_router_005_src_channel,             --          .channel
			sink_data          => id_router_005_src_data,                --          .data
			sink_startofpacket => id_router_005_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_005_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_005_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_005_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_005_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_005_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_005_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_005_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_005_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_006 : component nios_system_rsp_xbar_demux_002
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_006_src_ready,               --      sink.ready
			sink_channel       => id_router_006_src_channel,             --          .channel
			sink_data          => id_router_006_src_data,                --          .data
			sink_startofpacket => id_router_006_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_006_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_006_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_006_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_006_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_006_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_006_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_006_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_006_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_007 : component nios_system_rsp_xbar_demux_002
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_007_src_ready,               --      sink.ready
			sink_channel       => id_router_007_src_channel,             --          .channel
			sink_data          => id_router_007_src_data,                --          .data
			sink_startofpacket => id_router_007_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_007_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_007_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_007_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_007_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_007_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_007_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_007_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_007_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_008 : component nios_system_rsp_xbar_demux_002
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_008_src_ready,               --      sink.ready
			sink_channel       => id_router_008_src_channel,             --          .channel
			sink_data          => id_router_008_src_data,                --          .data
			sink_startofpacket => id_router_008_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_008_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_008_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_008_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_008_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_008_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_008_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_008_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_008_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_009 : component nios_system_rsp_xbar_demux_002
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_009_src_ready,               --      sink.ready
			sink_channel       => id_router_009_src_channel,             --          .channel
			sink_data          => id_router_009_src_data,                --          .data
			sink_startofpacket => id_router_009_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_009_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_009_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_009_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_009_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_009_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_009_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_009_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_009_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_mux : component nios_system_rsp_xbar_mux
		port map (
			clk                 => clk_clk,                               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => rsp_xbar_mux_src_ready,                --       src.ready
			src_valid           => rsp_xbar_mux_src_valid,                --          .valid
			src_data            => rsp_xbar_mux_src_data,                 --          .data
			src_channel         => rsp_xbar_mux_src_channel,              --          .channel
			src_startofpacket   => rsp_xbar_mux_src_startofpacket,        --          .startofpacket
			src_endofpacket     => rsp_xbar_mux_src_endofpacket,          --          .endofpacket
			sink0_ready         => rsp_xbar_demux_src0_ready,             --     sink0.ready
			sink0_valid         => rsp_xbar_demux_src0_valid,             --          .valid
			sink0_channel       => rsp_xbar_demux_src0_channel,           --          .channel
			sink0_data          => rsp_xbar_demux_src0_data,              --          .data
			sink0_startofpacket => rsp_xbar_demux_src0_startofpacket,     --          .startofpacket
			sink0_endofpacket   => rsp_xbar_demux_src0_endofpacket,       --          .endofpacket
			sink1_ready         => rsp_xbar_demux_001_src0_ready,         --     sink1.ready
			sink1_valid         => rsp_xbar_demux_001_src0_valid,         --          .valid
			sink1_channel       => rsp_xbar_demux_001_src0_channel,       --          .channel
			sink1_data          => rsp_xbar_demux_001_src0_data,          --          .data
			sink1_startofpacket => rsp_xbar_demux_001_src0_startofpacket, --          .startofpacket
			sink1_endofpacket   => rsp_xbar_demux_001_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_mux_001 : component nios_system_rsp_xbar_mux_001
		port map (
			clk                 => clk_clk,                               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => rsp_xbar_mux_001_src_ready,            --       src.ready
			src_valid           => rsp_xbar_mux_001_src_valid,            --          .valid
			src_data            => rsp_xbar_mux_001_src_data,             --          .data
			src_channel         => rsp_xbar_mux_001_src_channel,          --          .channel
			src_startofpacket   => rsp_xbar_mux_001_src_startofpacket,    --          .startofpacket
			src_endofpacket     => rsp_xbar_mux_001_src_endofpacket,      --          .endofpacket
			sink0_ready         => rsp_xbar_demux_src1_ready,             --     sink0.ready
			sink0_valid         => rsp_xbar_demux_src1_valid,             --          .valid
			sink0_channel       => rsp_xbar_demux_src1_channel,           --          .channel
			sink0_data          => rsp_xbar_demux_src1_data,              --          .data
			sink0_startofpacket => rsp_xbar_demux_src1_startofpacket,     --          .startofpacket
			sink0_endofpacket   => rsp_xbar_demux_src1_endofpacket,       --          .endofpacket
			sink1_ready         => rsp_xbar_demux_001_src1_ready,         --     sink1.ready
			sink1_valid         => rsp_xbar_demux_001_src1_valid,         --          .valid
			sink1_channel       => rsp_xbar_demux_001_src1_channel,       --          .channel
			sink1_data          => rsp_xbar_demux_001_src1_data,          --          .data
			sink1_startofpacket => rsp_xbar_demux_001_src1_startofpacket, --          .startofpacket
			sink1_endofpacket   => rsp_xbar_demux_001_src1_endofpacket,   --          .endofpacket
			sink2_ready         => rsp_xbar_demux_002_src0_ready,         --     sink2.ready
			sink2_valid         => rsp_xbar_demux_002_src0_valid,         --          .valid
			sink2_channel       => rsp_xbar_demux_002_src0_channel,       --          .channel
			sink2_data          => rsp_xbar_demux_002_src0_data,          --          .data
			sink2_startofpacket => rsp_xbar_demux_002_src0_startofpacket, --          .startofpacket
			sink2_endofpacket   => rsp_xbar_demux_002_src0_endofpacket,   --          .endofpacket
			sink3_ready         => rsp_xbar_demux_003_src0_ready,         --     sink3.ready
			sink3_valid         => rsp_xbar_demux_003_src0_valid,         --          .valid
			sink3_channel       => rsp_xbar_demux_003_src0_channel,       --          .channel
			sink3_data          => rsp_xbar_demux_003_src0_data,          --          .data
			sink3_startofpacket => rsp_xbar_demux_003_src0_startofpacket, --          .startofpacket
			sink3_endofpacket   => rsp_xbar_demux_003_src0_endofpacket,   --          .endofpacket
			sink4_ready         => rsp_xbar_demux_004_src0_ready,         --     sink4.ready
			sink4_valid         => rsp_xbar_demux_004_src0_valid,         --          .valid
			sink4_channel       => rsp_xbar_demux_004_src0_channel,       --          .channel
			sink4_data          => rsp_xbar_demux_004_src0_data,          --          .data
			sink4_startofpacket => rsp_xbar_demux_004_src0_startofpacket, --          .startofpacket
			sink4_endofpacket   => rsp_xbar_demux_004_src0_endofpacket,   --          .endofpacket
			sink5_ready         => rsp_xbar_demux_005_src0_ready,         --     sink5.ready
			sink5_valid         => rsp_xbar_demux_005_src0_valid,         --          .valid
			sink5_channel       => rsp_xbar_demux_005_src0_channel,       --          .channel
			sink5_data          => rsp_xbar_demux_005_src0_data,          --          .data
			sink5_startofpacket => rsp_xbar_demux_005_src0_startofpacket, --          .startofpacket
			sink5_endofpacket   => rsp_xbar_demux_005_src0_endofpacket,   --          .endofpacket
			sink6_ready         => rsp_xbar_demux_006_src0_ready,         --     sink6.ready
			sink6_valid         => rsp_xbar_demux_006_src0_valid,         --          .valid
			sink6_channel       => rsp_xbar_demux_006_src0_channel,       --          .channel
			sink6_data          => rsp_xbar_demux_006_src0_data,          --          .data
			sink6_startofpacket => rsp_xbar_demux_006_src0_startofpacket, --          .startofpacket
			sink6_endofpacket   => rsp_xbar_demux_006_src0_endofpacket,   --          .endofpacket
			sink7_ready         => rsp_xbar_demux_007_src0_ready,         --     sink7.ready
			sink7_valid         => rsp_xbar_demux_007_src0_valid,         --          .valid
			sink7_channel       => rsp_xbar_demux_007_src0_channel,       --          .channel
			sink7_data          => rsp_xbar_demux_007_src0_data,          --          .data
			sink7_startofpacket => rsp_xbar_demux_007_src0_startofpacket, --          .startofpacket
			sink7_endofpacket   => rsp_xbar_demux_007_src0_endofpacket,   --          .endofpacket
			sink8_ready         => rsp_xbar_demux_008_src0_ready,         --     sink8.ready
			sink8_valid         => rsp_xbar_demux_008_src0_valid,         --          .valid
			sink8_channel       => rsp_xbar_demux_008_src0_channel,       --          .channel
			sink8_data          => rsp_xbar_demux_008_src0_data,          --          .data
			sink8_startofpacket => rsp_xbar_demux_008_src0_startofpacket, --          .startofpacket
			sink8_endofpacket   => rsp_xbar_demux_008_src0_endofpacket,   --          .endofpacket
			sink9_ready         => rsp_xbar_demux_009_src0_ready,         --     sink9.ready
			sink9_valid         => rsp_xbar_demux_009_src0_valid,         --          .valid
			sink9_channel       => rsp_xbar_demux_009_src0_channel,       --          .channel
			sink9_data          => rsp_xbar_demux_009_src0_data,          --          .data
			sink9_startofpacket => rsp_xbar_demux_009_src0_startofpacket, --          .startofpacket
			sink9_endofpacket   => rsp_xbar_demux_009_src0_endofpacket    --          .endofpacket
		);

	irq_mapper : component nios_system_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,       -- receiver2.irq
			sender_irq    => nios2_qsys_0_d_irq_irq          --    sender.irq
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write_ports_inv <= not jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write;

	jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read_ports_inv <= not jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read;

	timer_0_s1_translator_avalon_anti_slave_0_write_ports_inv <= not timer_0_s1_translator_avalon_anti_slave_0_write;

	pio_0_s1_translator_avalon_anti_slave_0_write_ports_inv <= not pio_0_s1_translator_avalon_anti_slave_0_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of nios_system
