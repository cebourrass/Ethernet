configuration counter_conf of counter_entity is
  for counter_arc
  end for;  
end configuration counter_conf;