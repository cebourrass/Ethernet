configuration ticks_generator_conf of ticks_generator_entity is
  -- use work.counter_comp.all;
  for ticks_generator_arc_1
    for all : counter
       -- use configuration work.counter_conf;
    end for;
  end for;
end configuration ticks_generator_conf;